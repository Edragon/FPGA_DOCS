��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`nE`{`��u*���:�Pc5��W�^�s8�Q�\����y�X���eq�ym`�C�3�'ض �lM��~.B�D�@B.�V�]��#������BW�.��x��#����H��p@<��h�-�� ���䣥$�Jamu�_d�۫�/Q&lWm4|��āg/B���`T��_5�@k��M� �!��*^A*�J���w����綊�I�Ⱥ��O�|��/�i�����n�߆��!�c�n��+�-��<�k��$4�PUܓ��D<0^�� ���Vq]p�E�X�H#�Ķ6d�Vj;��>b�D�A_R�.�R[�{#�as�RLg�ё���LKƲ���|x�/6U��D4� ����Q���Cfk 8�����]1e����]����⩎� �Z|�}�G�8���u���_��(��F�r��v�[�ܝ�[�vT1seǝ����Xz�e�A��W,:�0DXkb�������Rv�ok ��c��s5��m�ux�>������\�����+)�.r���-��Z�@��=�o�e�'e$�c�r��̮�_V����;M�����w7�UX�i�u�tj( ��歨V�C\�a����X#r,���9���RC�P��Q���3� ��[�S�����T�MyNՌϫ�q��"_���!����pW{aKռq�@�\#�cPm�x����ev��~�i3R�$��-۳k��W��<�4M%�n���~�C�V##����'�wK�B�&��`!i���v׳2�����@����[�uܲQm���\�-�}��e��m�W.<�6���z����o�nv&�?=|n����/��3Ȼ�M�$@�|��$��lD����1Y��|��
؀w�Ůk���c.������,����Fw���x�}F]������mb��55�>a� nI�sc"U$��)-"�!vã�R<�7� ������Q�J����&��7�&����H5趴B�����H˫h��U�f��::�����.�[�gn2ɴ�n�l���X��J�uJ�~�3����	�����z9�,��f&C��sM��d�So�H06~�oǸ��E�����7ʣ�~ �C{�m^���D����<\wN�p��s�&�Bv8]���ƋD��[�M:�UT�����Z�.c'���P A�qB�|G�i
����N��	�=��!��M�k�0��Y�
:1w�xƁ�qc��tT�qD q㫛�P�*�mm�6�`��8oiT�J(�9 *����dkW�Av!��`��?+�:�d̍oH�q(	��7�&^X�����9�h_��v>��i�9qu�q��/��yT�oeq�¬��[).$����5���7�Hcw��4o�&�+�-:��!C�[Z��u����%}�`G*�熏Vi�wQ#ץȵ�:�0�����Z�؝Ϝ��_H j�s_0c!�����J�-�-��oj�cƝ?k����Mb���}�E3��C���{�{���8���ҡ,/�`�PF�E��� �s���@J!_eσ<5?fa�6�@O���lE���%��_ϡ���O�p�`~{`�D;���~}vGv����li���@�C"�N�S觴��*.-]�9�u��jTiA�������Wz3^�(΃w��HܝA&�����7�	�9� )د�:d�B��֕�R���/l�qE�H�h����E�.�ޮ��X
"�.�r���7J�Ӡ;gq�qn����O���3�+�M��v���Y�"e-�#�w����?����CE��X
mo˔����:֮��('�И06m���CΉAI�r�-o%uY8Kh��5i\�ׂp��3{E�)[���	���~�R�������8�I*�.�E)g�nQtJ��K��/	R�:?�ऊL]p�t�Ri`�>�n#J��������
�I#�4 ��h��&���R�?��G�b*|�:~��X{,M�W(�;��t��þH,��DO��2�LK��3��$�3��2�JMw�uKU[!�}�	>(�0D;�Jn����dDӡ���*iw6,j�I։��@+M�Z_?�ȴo��RBEH8�I����""��6����J���νR56�ټ��]�D��(\U�H|�RAc��%o��"��`��M �8��o�+_b���W8^��}����/U� ����L;PIDH���~Cs!cĵ�� L0Gu��������N�q�M�@�~��+�/;j�M2�{���ʀ�n��4�r�B2��ɢ����'� \����+�凧��}�`��[N4�0}�����0��O����"{�=�|I��*+�^,J�X_B�SYeS;�V����RKO�o>C��c�:_��!G�M��DMFv�̩a*�j�M���{=r�Tע��(�	�g���t
clKh��f����e�8�����Kb����.��5�[�2;G&��`bڧ�\{�)�K	��P�� ]�&��x���h#�gI)���r5��*4\����`�EeqR:G��[�w�`6�Z˵(*c�J���[PU�/U���<i�\@ƾ�0��Z���G�q���ĩ~q����q�»:-Q.M��+oc2Air�cV��D�FE�,}��3q�85ϝ$��p7�G�V�}9)�v��y�~�0G	�Խ��nZ���b���ΠN~�YC����ͳ�Wn"��'�S�K�9��A	/�Q����h����3C�GG�l�j�@w`L���1w2MaS&�P0dy��@&�>�2";��K�n���8	��� ���z<�W'��x�s�p[!�����5�e����z�
H���En^�s���l����H���bj���s|�.�٥q�4���g���z[i�	�vÄٔ�ԲM[;t��q��=�㘉꽚E�#�̲;	�6�;h�ߛ厜`�y(�+hU���k�����`�43�m޸*�b���*�2����"O�~�ӧ���3�$ B?�:�`�����-�~#Ӈ�<3�ʞ�{����%���6�jIԈ͉T�9� �KH���$��y	?.q^��w��[a�j��T�tC�Q�V��?;&���Ѹ�7���܆W%f+M�1hF�����΂��S7�i+vK���#�����u$!��&���AȲ{Γg���ne��'����$��=�>aGc��|��!o�5g=�����tv�'��s���I�Ϩ�W
cЋ��G�]g�ma+t�,���C��ֲX��R�ς���TSD�ݥY�!�v?ٯ��Vz###}��|	.d"�&46قe$�y=��;>�!;���!��B�Yy�Hd#�/�?}kz���E ��<�"�&t^�K��odz#C�u��ĝG�	���Pd��4��Y� T�����*�3[Jaī.�F�^Q�lJF�����֦��:�����\]%����,���j�P�̡�P�n�q�+f`���H���ͼ�9���jA�2���Б^c�S��q =�A��[��m�[��[X�?a4[F��P��LIu��;d@;���D� �Ź�R{�.�{h��[ �NHr;��u;��D�@�&�����#����c�9خ�4���D^}��y��.S��8p���y���%U�&j�D��#Cn����=�(/��ɛŜ˂����72�<���8K�8N|� \��w����@�^�oy��p:�7O��]�ge����/Q|���/$��ևd����l��6&l�Q[I�1�p��7/����g*^��۶q"^�C������,�n��T*�>r���\�ߏG嫙�LZ��	DO���x�m�|�@�N��v�g�~;6�1�w��?=I����`n��ƒB�/7i���ǫ9o��eX��&[I2���sMa�-��"�N���kg�	yϮ��>6�)O���ax���v�{1)nK*6e��rC	��/�u��'b�ݟ���f�����xh��V�j��T�bj"���b��Ŧ�[����)S[�`��.����w��K��"P����J#?�"��E\�_c��_��o�`��IC0�C?�Z�h���
�*r	�ɯ�t�&��2HQ:�!#1:����R�s4�J���,�C�W�5��WJ�����Gb}U�qm�]l2D����(>�fR�l#�ÞKKW<H�%���iO�M/�;֗$�j�RG��<�d�W�gm�=�"�����=����|W �~���tx��M0��v蔉�t�n���E�/�l���
��8uG#~&5���F��3��\�qs���>��~5��wD	��f���uXR�D8UE��m��{�VL)qNL9o@[���9��)��ޅe1��"~K�&�-�a Xx�ӕ���Xi}MH7����9q՘��I�xq1V*�u��4��\J�,\0t�6��A��(�=W�XRZzq%;�'�
4�4zLB� .oYdrE�;�q�̅T~H���/i���j��^�"3�3��;^�=�(j��g~��^Y��pẊ��U�,��`�����]r	�&Xy��C�tW�$�8p(Fe�_ ��-pLF���8nB^��s���4���4TÌGϔ���FU+� 4�w�1QD����БkD�,�,9_��%[Y���$Sމ�i����U�hhH^)H�[s��0(]�1W���$:����cs@d��):���ATv�l�u�������w
�����v!�ԥ�pv����J��3��V,���Â,ى<�|Q��RK�[��/�/����in�!�L�|�;1�6�rf���q:'����~���DI��L����qy����A	�3,��Q؊��5E�� �g��~�q�"��vK�@l���-�D9���7�-~F�������b.��_=��ӳ����~Ė��:_x�p�ث���}�X4��3��}s����9�̇u��O�b(f������wb�v�l�V/�-|m��Y��s2��>�	½�Z��7iÁñ/S�4�͋q7$;�7M���̕�� ��3g3��"	�F@3F���l����֮���u�>^�1A�s��T�sֺ4}��C���ơu���D)I˙�h����������-�e�%���M��"A���1�3ͷUUf���2*�_}�W��L��|jRĪ��4o���5�\�]
��/c�'W�S�$�����!a`8��;l�<��^bzsv�p�#m�?���7Cx�9]T�d�jb�K�,ױ��A�F�e%�Vc�pyx2��W��H��ki��Z.��K�����1.���[����g�@!z��|�w�bk����G�TY�%����\�8�����J�R��u�y8�T��ñ:�4
֕��
g⼋{�*�[ۉto���{N�+��9�A���&��v�c�f�Y5�"��B�|�a��c�5N/q�}����t�����q�]G����I��.���l5��V�%�N�2t%w�~�p�O]�%Q��E��e%��{��-�{�ߘ�}߯k�HU�A�~�0̬��[ ��Z6ug*�M��"���OD�l������rI�e=<��I&�5�2�N���
�;�cR--��Gd�6kW=Ov�m�I���C�bɂ�����%�;��>���<@_����$f>��+b��M�@�Ҕ\��n$��*@J"�	�|�|�}	�����0!]���xª�W���Fdt3�~g�J?�(��U6�o���I�V��d7'0x%��vͯ"ݭ3��t;rO�W������sb��ﳙ&��1	������]Qv��"����%����0����c��*J@�l -!8
�ZX��ZR��>�%9}0~F ����{b��mk�JMc#��=�ɰ�0uF�]⁗AQ���K������I%)J )����SGn���w1ʐdI�71�;����N����VSK�����Hmq�9��W���AX�x��;R��{9Ľ+���h�:�9r2�tV�c�U�E�4q]�Xu��O��hʀ��I�D��ij���њLS6��L�u�q�r>�M����ۦ��U�i?oR4���:��<h^��g���z`�:Y��%�AO���Q�2�w�U�3�JP���K��6��uV�	tFj#��i�
c�iHق�!�����g����¾8:�{Di\)����f��݌ ������m9+8�}�7�Gb��i���m��۵�h���Ք	>���Px2������p���!\��n��_J�j��^9���͟�g�1�Cg�G!��|p��,��`��ל����&�CJT�T�?-�w�ɐ�����ʺ�([�]��������c���9���lrj�X����]p��ȍ0y5�]�qC�Z*l�1/�����Ȁ�`�GmB��c�Ix�Q��DW��'�:K�c�3�����lLD����.W�8}Zkd(��sYέ].*���CX&yFU�9�8�UL�����4���j���V�I��@�sԀ��4���f*\҈qT���|��
��h���Ph�\(Rl������j��k�
��	�"�^x
�w}��B_�)|�\���MT�J.�ķd�4ˋAt�_wDS���R�"p��:�B01�3��� �L�����K�\#��ߪq�ǜ(/ы��#��Ւf��q�9J\B��v�\r��:���a\�Q�����qF����d�R&i��>)�mӵ���$��ܟ�=0W�u��Iٞ�V�礶�� M:�Xdv����S^�B�BN�f=�ޥjKU�D�+�����p�p�p؉�
�,N�x"�_>j�+y�b��5W��zi���&�����20Vc�R�����N���:ܿ�[�[݋��<��|�8�}�-���z	v�t�裥���gqą�I� �`Uo�9�|[4�/a��'O�����	k�a'�Ӏ[}ȼ�$iL�yw-���i0f�m�ƴ�I�׳Ōr�|�q����"���>�J�2��YFRȯ�b�`|8]�%yQ���Ӵ��!*8�oG�����#u��q5A�Y���Hbn���G�W�um��)�#>�Ns֠��o���(|��j[$6�<:�6��PF�׃)7�k~�}Xl5�Ew���3g��_ੰ����e�]x��AJb��(5v��Q)���O�=��l?S��W�}�d��`�~R��؎��H��Б���-\w����t��Ș�?� '��>�.���m��!$��uW�r��z���e��oύ��"eeZ�q7��u�c�9E*�0=�'�h `:��vaI'���Ș��8Y4K4��V<:���v�$c0���,p��e�kw&;qy:�>e<�~}!�7����6�$��-�n��Rl�o�D!����pp�˧^HaS�����o��8�z��P*M�x�	N�,��z8}������89�7�:k\Y�f&f��9�IyB���D��XJ�V��ĺ&�&e��l�e=�Q,��Ӯ��d�-P��������/����hCH�x�\ �~���S��ٴ�S�L�gd2K��x����~�!H�>B�AXv��?�t�*V���v�p��	c�&���#(�1΁Ñڕ3RcC���/�6�3#���������:K��H"��|ۋ��	%��� S�ge�^��pj���F־�S�5�չ���HF��t�#}�آx�*�Y���9�0ֱm�戔2�N������ݳ+�L�>.)Q��5F��-K�8�:S�V�j��*�U�n�cMX�����?�B?���bX���Q'���C\x��/l<�N�� �;M#W�ۈ`BXm��Y�>��^�簹�z	(�L���|0xfK@WpkL���wL��U�t���M]�[䝀���Z?���zh������_؇�;�yR�ȥ-�>}��O�!հ	�H�(���s!Wb�����j�s���5����=cC�a"&��
4�������giY�}-��y�%�7@O5XA_���ȁU�9%�%����E�.g1'!����x�*z���g� ��8�?e��_8�U��@�P���~&�U[�Zd��Ȇ��-r��]���g+G�0��ZUq����̒j��>t�m�]�Ucb�DQ=d�	��G�%G�$rդ�fƠ�꠫��6�,`��� �\R�f+�d����=>�c
�A�Ղ�Ң����X���u��y��Q}<�5-l�֚o��7G����y�r��3-J���;�",�I:��L��㦳+�螤�5��	=n��[���4�=��L��ZSĲ̈dAΈ?����=b_��8y��{\Qh��Z:���-�a� P�P^��0����B*"����ک�Fs )h�]����S���>�Q�N��c�k�~B���)Ĥ1wj�vp��Ҳ;�B�H����U��B�<s�JTL��ET*Ϗܛ��	mq������.�2p�Z�N]����ӁL���5�l�4FY&�젋�%��)��G���f�3h� ���َ��W�u��Z�gx2,�P��&��2[�	�u�R��ȡ*��O֧�'������?c>�+�/�̥4��`̔����g�K.xa����[��=s;'�L�C8xK'*E7�1�r�Ǭ&Q*:*�)*� ?�ޛ���i�"K�4��\[H�.\+���ⴹ�V���3)jGo�!9��Z��Bx���ucXZ'#�ۨ��O[QaE��ԈQ���%�%X�]$��q���F��(v�ݥ��ཻV5:}X�@��H�~6-Ⱥ�$���-�x��Z�pl�����s��s~�r��R�$�Ik�V�p�ί8�]eDDt"#I]�@��J�yalL��#�:��[._X3>@6��l��F��9�I<Q.��q����~=�{aNھt�N,͢n�?RҼi�����$�ǄA�/^���T[]`�K�]�ܠ�G�4E�}�Q(�C��H,F���tu�5Cgݮܞa�d��V�Dm&��^�f���D�G�n��'��_��Fj�v*1 &�Q��(������ˀ�HS�mO��CD����_l�8Ǯ��C�\�A�KH����5k-˶�>���0��6^Bn��Z]!DX-�ǉ*TJp�{��G�5�j�}�[`I�lyl%�e��-���z��FV���_&�6�!t�{Pn``H������3/�?���Hu�P';yw:W>�|��F���:�qj�)B�Y��ٿ�s8fvo+YAY�wtsro�_�&��D���
��5�Wˁ�˓� v_���a�a��,����];!d����$�:TL�TT�P���ep>NGT� aV�,R:��Gq^��&�9��[L����Θ;P`��o���Ȯ�%��c[Rem$M/�{
Ap����L:������=�����f(k2E�W��u+b�Z+1Z�ݡJL �{��8�g����5��H5:�l�s#�3�:,g��7l<'���r	���'�F�2䖑B1V�t���̈:��;V��$�/�,���]�<ݼ�����֮���L�NU�~����^C��g7������C���K9+���)>mS�Ltݲ��h�Ay^4z� 	���x�z��NX�|k+��(J�����P:�a��}G���b��N\�OY�X�e����H3f�Y��/�,�����Ҡ���vW��,Cj�<**�﯌p��4kP��p���z��+�	 3R�4�&�Oq�r��gW:��l��WP]�H���$�fY�?Jw�(�U�ɔ&�����3����tX��B㳬0H
����p���\�ai6
�%�r�*9T9���?���I��l��/�)���3����pJY��w����,3�k��`Ҧ>`!~��X����캭ߔ8X��Sx;�O+6�S��:����-)����d��c�-bN���u5m�.�@S��|�u��$%;H����_b�ѷD@�b��T"��X#e�y��������i5]��>��K��eb52m[�x���<B������/�[�vr�	�,(y��v�>d���X�햔��A��4�ȋ���j�_�:'�u�:]~��ݘf�J"��fm����~��� �CYVa.cs���M*3�Sn�U����'�������;�9M��
A�V�2
+aE�3�}:���m�3:>ґ�A����U�)��{O��A� ��;�_ڴ�����j��f0�A!��Zu�V�	q:�N�9��\c�&�6����,�B��*9�����6�"��C����O�c��S��,N>����'}1xT�LK��_<�O�j:�vĲ�)Fב[�����m��UN�^�'�	���c���zZ�����)-ˌF�q��"ZuB�L��ܤ�l�7�OO��d���R��I���fă���,��"���0�����!`����[^6�R}k�6S�dq�&�X�`I(��64�]6Ȟ���Z	P}�0؉���:�؃����n~v: cj��J��@,�e���	GQ\���Z��L�Q��Dda��������{Y��o/)Q&�y�p�>�i(��;�j<��Zf7�I�K;��N%� ��'�`��O�ZeOK�ä��2gYoG/�̑�*^e"\O#��y�l�(�VFz�d]��m�q��ɓV�8�A��w�U��ߟ��"�u�)�hݝ�pqi��t��݇�I�������Ⳓ*�2���w������������!�־o'�WA��HE����:p �D=���i��.V��1��䣢�l�����!Q����2*(_<iy<����,����X��,��g�I���AjQɰ5#
�PP��F(�]K���r>�fNCy��X!�q�B%LI�j4�<��>WO���Hl� �Ki���i��#փ�T���ITi���;-��(��39g�E��؜�_^�ߥ`����t�2O�rϑG�]�l��2ȷ#�H�fn+��)-� �YC@��^A�T���zNb"R �$s����B�_+1��+@7��s'��v��0m�����)��|��y�����ԫk�$e�U�$\|�&��@����I[\�R����A����֋j�@�a��"L,5i��oD ����G��

=����@H����n��ڇ&37Pa�B-�G'������Sb�H�[�-�$�u�����}^ ~����-X,*۟��c�Z�1L���Rk���֦��8R��?�4��@��'��\�p�Un�vB�~L:N��b�ɵ��>4�E�f��Al���}_d0��Q��c71�SE�\�|-����'��Ĵ��6��[|�z�w�澄`qR��[�*k����F���`��Y�3��	�I�R8Ӌ#[p�����e�GU ��^�5J-��@�s�� �+6�C�(6>슕�4��3D��ٲJ������2C���Qɱڴ4������O/���	��	,�2���|j����)�'%��\{��h
�����&2�H}v�_m(y�8DdhSҖW�ZHj*�I��=�+�5߸2� -]�Љ
�o7�M ���n�>­�lǓk�x��'j����%�<�j����������o�W+~23��p�̼#33}�1�{��<��-�"��^���kJr�y�j�'K_/'Ү��,�Kҡ50N��0�b��e����A��4��z%����̥�a�F<�;�o�4'����k7K�Ρ
u��#�O��ޝ�N�#+\.7pJDi 
�F�jy�Kq�pF_�x��M"�P������n�b^*L&�z��`{>�zI�x�yx�[�%>rĠ��3R^w�3�yl~�܅��zT)9�%F�A�>p`��i��&��*���h���y3�P"�d�N �k'�5<ax�.Z�(�3����6�7�����o-��T�'<�rr�ڿq����Nq
�`r����E���Tڧ%*���/�{ɍ��~_Vq�i�i��E�r��)7�so����R� cL㑓���Rc��j�g+��nP��'���G� e<�$�|�����ٚ��Gɷ��b9`���5�8�y8�tr`;���|;7{�[_v��|�ee���g߃�JDI"{��7���W�l�� ���4��V�C��y�,�#_��M�wR�)��x='���M�1��Y�uG������$]����{Q���n�X�ǂFh!�-@p[W���|�'N��x����7>gT}&=f<A�H*!`m�N@۫���i�>|�����c��.�c��&�q�߂�o�8�;�_��hJS�8^��(����+(����"�hÌ��ª=1��S卿l�/��Im����r-mf75�Sf��,�R;1�>��"K/��T��<�쓈�=p���s<+Գղ����$'/�'�H�l{;��*��Ie�_���$�Jچ�o�=:UkΝG��oB�?��Ƽ[����I�yN";�:��n���;�|t8��&�)O^�ѷT�07�^��qd�b��P��� �J\
����$���o�Z	Ik��\���"<)�㪲 ^ �:��B.+<!��((�R^ވD�\��{0<�,��p쥂c@4A���2�|���� ^C��v�3<���u��y�=�3�?3����!�W��>��>,%�����e���9�ٚ��=�R@�w%y�Kl*��6�J�񬔵��8m�`P�	��B�Q�b2"	�t]�7�ޖ3���<�@��|Y~���������	ZH�H=��\��� ��Z��yē���7����?�+��[)��t�yT
�3^�s݊w������6�@�����;By�voѰa�W�M�e����,��%�w�������\yP0�)���gx�^jA��usS=z��������?C�Ei�X�C�\th�f&!�Y%,F)���Z ��f<*|t���g����^��n���y4Zù$��><�����F�o���s�\�+�$I��L'�l��lB����yLgG�ybę0;�9�`}{'h8K����0i�`��#5.�S�%���2�/��i-�i,vѰ5�[x�I7�����4�R[��Í�����-P|��E����6�]�b�w.�șJN�&���� ��GX�j6���)� �Q�[{���)���0�����wHy���#uC/Swe�CfMr7D,�ܢ���Mǵ�~A�/炥��#<�1��V�L���7l@�L�>��}�����8k�:0�Qǥpw��p�^X�__`���J��+�T�𽃋Q݈ͧRܥ�8����F���#��"E}:"�[��� �;�#qHa��O|u�mEԠj~��,��{�3����Mp�\���]!�N�0�ɕ���L���6~�PB4���%�m[��D7���ӿ��$YWr ��� >K���r<3cV���Y��H�����9����{���l����\{3|-�F�MOE�@f���uO��/ո�!"?X��ۻ�w���ڤXڤt�3�H�;�&p��Q_u��C��7�7��ҙV�r������r'˥A�a~UF6����#��6�>
W:�0$��ۆ�M�Q�B�� و�k��@�9��ɜ$xD��n�����A�~�>�	5:�~�Ȼ���������%0%E��[�D���R؊u_��2i1�8��goA0��N�X�ޟ��A�k��R�5�1ݥ+o����� i����o[F�1;��V��V�;�6|�|�.-�-㪚n�\�b�ڲa�Z@ȟs#��"Uԗ������~��t�>�^�+3 ��Y,f�)��dЉ��9�&Y�Azn�$n9em��c&�\�vkQ�#��;*� ��C[ZѾ:?��'i3u�k�Ol����v�`R��q9Y����������>�O*h��m%Y�����[D7�˶ֹ���x�o���$zR�g���DG�g�e ������ͻ?�����Z )�@kh䅛?�\�-֡�Y���\GD���)K]��{ 2M2�u�,;�W3Ƅ3t�����3D���r�&�8z'8��@D3�~�uL��aN�N`�8�¬
yy��_��,4#Z�/挶#Z!m�a&$�$�Ή��K?���:�T<���V�Xw�%rg.;�D�Wʻ�/�}�`KR& &`O��QUy~>%��.�L�P�?i���6/���_T*Ko
�����~�^��R���Y����Rcj���[�G��Q�k�3����������;���@]�s��-��9®�j�P�ՒAI����	V9�e�<����4�#p�pk�8�]a�0���Ƞ�P�U9&�;������>���lZX6����:�p��<Û�h��`x:8F�H������I4�PEP� C�u�ۺ,^��2H�V��Y��P�E2I�Ɉ8 �~-�"�UW��Y�"�Uk����Nb��*^6|�b��{�_��w-�&`�J�XH�u�z?X`���Ɛb��J�[i?��Q+�&I'H��0��"p<LE��|0} �^�˭Ш2�i*�Ib���1ӂ��Q��ҹ+yÁlM���s�h^S�9z,K�q^��Bg�EY�*7;��pm�8"k����������,~��ַY-�%D�j�Q	b�����zKђZ�/ػ�)'ߧ� _�/�ڼ�M�C����K8o!E(�0�p��S��n^���%���p���io��WBN��ߟ����EP���"�B[Ii�9r�zU����O�� r�h�n:��9jC��:@n&"�$��Yib���w�Tv+>t�ٕ���쾐]E"�j,�QU���|B����!h�|7��ut���7ʊ|�n%lCҙ��|�N�v�6����o6/����{�����(��ޏ@dE:3E�Ӑ}K��%�|e(�/ݯ�`_W��F���z,RGez��i]��c�b��܌�:ȝ�1�1
k=m�#g˭����ނN�H~}2
*��q_U}eΓ��^��5��4(t=\��)zk�l��)_�"y��˼����{�Ӭ�d��{���H��a:*4�rv������v����9O������S�;)sBŊO$�o�%;
Eb�L����#@=]�?)�^���]2p�Rg��5������:�H*�)8�`d.߫1�Oi��V�AH��o93�'1�_ġ��u��K�X��7[_J�{n碀���a_,F��mc�t�p��$֒}���Z�g�`��iS�|��_ ۾����2��b��z!�0�m�G��X�= �>���T`��Y�S,c�! )Q����+@7�;���
5�#�	^�8\�O��F3���0�n�k���� �|��z������~���7��ύ�i�}��o�A�}�9>n:���P��+M!�dQ�g�ց���bb��6:ޚ8ea�;qO����������K��b�#i2T]ǆ�a.� 8���/����<�jS��`���j���DF�~hl�Rz�Ca}�"�p~ͷ"�M��������/�oצ�@�u���uݍ�.�������>[z�v�S�,��}�AD%�N��KTG<q
�
0�!�|��>ꢠ%\�[͓�/Λ���&��{dM��+����>��k6�˧�ε��ؠ1�o��Q�NND'
;��9�4H��`�@��9`<g.���x���,g�w�0K��Μ�Ɏ~!��9���Ss �!`�t�[�S���'��%z�´�7,�J����
��y�uX���1eX2z�����[jn�VH���Mf�~�T�]����K}zԏ�q�N}��.%Q\�H�~^�N���4� [S���V����Tc~����>���R8?��	��|7S�I^b��D	��!>��<���~D���#�M�B�Uƒ�� ����$�2 ?�4�p�t��U��;Oˢ�T+��e�[y��#m��F*ʖ݃P�s� ��a��f\a����0p�`w���[a�g��S�
��������3&u�3����V�A�������u����}��شŋ�f=�RvB|[��0H⡁�HvQ��*y.�|'?�v�NB��w�g6%��n���z�v�J����l���T��2>>�Y�&��$LM!L�6�K���o8�\x8��w��x�ր��;��cx��GVn�̃��>��P#:����-)St�}���R�Qs�����vX=U�e4K '-zz�۲݅�!�����MT{+�o�T0��3c�$7����#\��n�(iq���\�1&��+$�@�H�Ƀ3=R��Cc��qU�C7/Ga�t�v|� �3�U�T�YL�o��=/l	����w�pHut_�?��T7m]0qI�	넬�~҆�y��-
� 3R�omp)�''r����Yb{��7-� 6~T��)�-�B������uL��1��"j' L�5�3���C�����Ƨ���^��V�˄+��5��A� fZ�
W!�1�&�$y��$G�]dV>EQ���f�@�&>>�U�^�aY��}�C�>���P�c��#��\�d:������됭 ̚Cno�V�ӧ�E��̎Z��
��y�����L��Vƺ�������o��.ǻ뾌$G�U�����9X�=�L�j��ɑ�#���X���v�@�9�Sl�nh�Aa$���i2 fx��@7�)���a�v�`08�)��K#�t���T���VTXy��C�_��]D������X�c8冨
��)ஃ=f��a3���� ��t2ԯ�v��0洁�C�dʓ+���e��~��£��n��lsd=���DPSK:�zx��q �k]4 ���q��;'�r�IR�c?�߲N\:�G;���Z���+i���=ԋ�ۼ��+9��S��2b
�#�H;��UU�BgDį���|�R�))J>x�-����2�*�c�6�=-PA7�H���^{v)'�7a���$�)oL��zJ��h����fAmc�1G�=�� m�z�|Ό`To���뀪S�k�U:�ʨyQ�V^�5�mž�Q�e"�K���M�Z؟	��Z�����v�	h��mm>J�/bZ	�sW���(Z�5?�eݾs���eD�gp
�^�Ψ����/Xj���v,k�a���WTʨ�rI�_�09�)��g��*[��=���hCG�"p+!m�MZn��J�]Y0�u���K�NW��#1-�/X��������E�李&o�l:����el��Ŋ��g��{��+@�0�}�/�}�!A�����S���R7Da:f�����˪`2�5�����"��L��cl'T3�p������ ���Ưh/E�4b�u�
%ʰ_.`j�rD:���8�� {���]���^tb��\��+	�7�����	{3��}ng��j����!��Ě�$��Am6д��ū��q������;b*�_�����ŧ�F������N���	~KW]-@g}���YP�V�=od�k�q��4�������Q�#n�c�jx�������6��l��O�?5Q?�j"7
�ܮ�F�ݼ\��3Sj�v�.ҠZ~T)�&�j�9�a�N��K��ǋ���@!�uU��aE�w`O�m�����e�(c����J�l��/kR*
��i���i�o0�xu$S� �!�-������p�������6�:�5]���Ϧ{i63D��Y��#[R>H�)Hd���f�����_����M�p	��VG;��1�G��͖�I-3d �$.���}�E� "��\��ˬ7t�+=A	�8+����쒸�����B��:x=N9<`fjZHy+�{��Lb�>|�	ְz��xP� 6$���L��O�NÙ��>Nil�p�AwK��:o����Vm%M�!�I�3���Pa��E��(��%�4[n:N���+��= ЁN��'�^k'� G�g�O���@�hE��������D��O�6�,n*��2՟�|m�ȣ����h���]@?�����u� yG�:;��z�<G�����]�pWm�W{��}l�svR�Akq,�74h�2���q�apzW{醹���Z[+U�N*�lF�?V�_δ���Ȧ�ݙ̨���}~WH���4�<���ֆ�?r��]�R�[�BϞ趵��9�`-�A��ݟ����zj����
���_Jn��E����1��9��;�	�ն��K]%��D�2�AOЃJThj�,��eVmHܮ���E?h�G�w?/��@��b��Hė������70�����جa>�	���g�U��h$;�(]�M/wqBc\��W"獌�(���"��e��:�;+(<�؄�ء4c��U��1~	O �]���Z��m��'����#�=�$�D�Y#�<8t��1<VFi?�Nc�>_��g3jċhӘ�����:Z��L���*���>Z�����b�5�jJ���]�����7vq�5�v�!Nk�o>0����2�����Lp�c��#����x^���=��F�ݒ)�\P��.�F�~��0��bLs�輫�w��������Q>��>p�4�!��gEWl��6�k�Lg��1�a�	_U&�V��H���#6�ƓL�o�n2������P\��������4�I_iM	��>����f-Wm)_���ir	�D����%��J-sk��6�JY{E�������:�Ũ�1��g�1A�37ir]m��]X��W9�4+�5���)�x�Eq����`��/�7���u4�ǾM	���h�q�`��T!Zԥ�PyxUZ��`KDp���-0��|ir�tb�S��֩�A0��#���M.�����w���!T9�DB6����α�����א��aZ��4������K/�k[�(Ԏ�ͣt
	���4N�N�}]b��-��pQ�"x����v�)��@W1��c�-_Ψ���P�p&�q�]���+�2"�UE:D=�r���"�x�.�z#Y�"B��<l8A���4J 
C����j/�N?��Z2��L^I1/���r3��#���q�3q#lV����#��PV�Nv��D/CH�e��k��^<R���2��e�ue]?�l�2O�$����iᆪ���\�ٖ��%���~j����H|
A�qb�/rUw Q�Ӎq�	��PY��ǡ��Hz�Y�?iǮ����D)����C��*	��!k�I��xzځC���CU�+U$u����'�a��b��_���[�:���X���=�1Z�e��D���V�O5X����.�bDSW�sb�ty�:vs���9Z�Z��D��p\,y[��el�� �O#ܵ�Ӈ?)~4_>�2�!�ȹ���P��6���)�����"Rr)�i�1����.m�:�d����S�
����@լWC]����*�s*F�ÆuF����V���#T��ew�Bnǯ0���Pi�������R�l��e�5!�ޤW�(\S��s�XW�[��poJ|Ϭ9@^T0�@ӧ]U}��dᑐM�s��Μ��N0��z��w���h��4v��uz�����Ce���<9^&���Q����<.,gIs=�4ߧ�ւEkx�!�`����P�F����>���`�*��
�Jng��z�2O@z��5�l�	��^�|`�69��_�M}�).��`�>�(�2������~��~8�vv��]�@�i�e���t��֐n ���0��C�Qy� ���!��3]��S��������u���<���~P���Bau���ٻ���N>����J���Й$�Tbr�l��嚥D3|��C�FJv<�vTOlNߗi��ڶ�ǽھ߸.Y}$m?�~�U�5�� ��n,�KŹ:2��͂iȏ�f�����ˬ��>��q+�Za�R�H��g@��
�5^2����M���L�{���v�7��"t� ��2�� ��;is[V$S~r4���f9����R[v��隍�2kq�U=����T� A��E7��^���\&S���D�T]`u�Qa4���V��n񧻈?/�?�J���OQ,��ͨ�^o���2�M�O�����M��l�_��@6�G	�	%�����e���k#�d����<�QmS�n��0���O���>f�k�m?�����w�,̌,��Ε�in��b2���c0W-�����0hع�3ի��S��/���;Ð�t-��� ES���Wn�7���SW�iL�'���H�f�������@!P�H��!��q�*�}�:ۨˎQ�Օ]���LGB�D�H�9��RA~X����<��d�p�V�ɬtǹ��Z�(Xko��'�e��xZ'N��E�p�V{����o'Ɖ��n U�����'��+U������X�_j��.YE��� �Y�
����@Dpqs ��|i�� ��9u�L�>fĝbr�^��л��MKM*���2���W�J[�B�|�ߤ�/P��뺋"���@�$�E����iו�YC�4)�qf�j�s��j:��z�����6����՗�x{��5�;hS}:��O�aE�n�Ҏw=N����R X
�AyG��p���m�Gh�d�r�Oz�K��W�Ω��+�F�Ƌ��,�_ii)\U�I�hX��)�/����T�B��;���,o�w�=�{}��@�\�њܑ�*��E�񷒊�܎�;SG�V�৬b����?"�eˢ߰H����$���*�j���r>��7<�=tERX�B�'8���\����Xd�.Ɋ?�H^���*찤,}�t�)����hЋ�G�XCҀ&I�Ŗ"����E6���O�r+�m<�y���U/�5��A����7�^�;ė�!�x�
v �G�5#�:
U��	�Tʧ8C�փuz�;t����q)�o>}\	M��vu�t�����+r�'�h(��!4��C�V���<8ZCdҔ�t�VLV��1�Z?�.��D�Բ� �[��A�	$��^JM�w����´�f3<�y�.3_:F{E��ɗN[��{��`#p��J_���OrL�l�Qt��$I�� '��X]
T�1�k��K�ɴ|��%�(Q<�r���}�H������xB@Y\��
R6E�����)�}�|��9L��̣�"�A*�8A����OH���)$�Q�P$��y�X�ax\�%rJ)+��վ���[��CPx�/�ZB�Tu���]����v~����n3Pl�Η�n4��,��E>ȗ���ME�?����N4�u��q�n(>��%�O�2��m������~�������]�)W���\���I}����y��s��]�1-:�3*��>����>T��� ńG�b���`�?\;��f�&+�'6�l^�%�uu�����_	9��Yk�"-���[0���*�@�I��&Xɤ�)uoG�@Z�#�-�@���e��p����n6"�؉l(C""3��5�ƹڲ�[;�?Ʒ�킄�W��
����u�"�L�J��pX���Jz�? ��.�{�o�!:�!�]�⁽��h�tr���Z>��}����M��}��߬Q�����z����E,�9vH�ICe^%��u��U�h�xo-K�:���d��̄���V���y��\V��r���KmN1w{Y�V�qw�`8�b� ��0W�����f�aU���'���Z�mB�dM�#`�"����\��$M_��4 N�X����V�I%n�s�Dg3�i^�.�x�,�}ktW���z�;����C}W��ؗV�+(+�k��c��8Z$|u]M<�ag� 7Q�P�`�٤�Ⱥy�ʵJ���i#$�?m���0{BM�5?l�"�C'Ɯj����vM����|S����F�5(5����-:�k�����Eܷ�X�/�̄*��6�/����7�q�������ʄ>�Ƴ�Ee�@�&a������h|�9~.(�;e譋ݹ�Q�2a�/C&1a� �{�&�Ţ�X�f��96Pw���D���i�t�@W�ێ�7r����!ѸQ
��j��B)�{Zr�z2�{%������oN.��G�y�_�Z�J����u����1X�MK��{��gZ���R�Q��<ۙ�R{��(?���Ta�Ӳ��⪞lLR���l��]�o�o�J6|K�f��jlL�=MK��j㙚�Ÿ��.莼n	��{7hzYRT"��Tm��d����b��
�<σ"w���]Lx򇍿��3�6 !����6��m[.���Q$�U����l!�E.�/x������S:K6	�:�'�Po���o��	�����81++17�O9����.�P�4.��n�uhKq�)�c�n�-��e�wP��Kf"I�
�Oj��IoW�\��!���<2�1���ؤ�����|;�g-o�}CN'�1rKKM=�M0�*j��L~_	�6�
_�_p���K��[%1��šC7RyX��������$Pk�H�0��?�f�۟�W�,��Cu��Ѡabt;/P6�l�*��.�cQwow(�,=� T���� .�z9�n8t^�[I�sy���NҾ_ �W-}��y�{��]�ൽr?�4�KjdS@��^7$Kw=��@n�5���)E���߸�������W�cp�ܼ�@����QQ����e�����ZĢ�"!�ϝDA8kxm.�x�D�ꭱD��7����i�~J:�ׇ��4����u��c�+��:�P�h�U!��c&9��U�`b����z��l�0[���2�1ܑ&����2N��6�<���
|� �����1N��T�6��q��H�j��T��W�AH�:a����8O�����Kbzh%�_��Q�s�;ʎ���RNko�
J��>���h��x>�VͽF��M��f~�����=Pm}�_�If��0b��]]+Y�RZw�#�G�UywJ&-o���g����A+���a:���C�򲯤,��\"�� !Nݞ���֕)^8��!��v9�O
�B�5_h�
�p1?:".ۢ�IP]�����a�ȸd����j�Z�9&Y���=�[��(8��2=��u�,�C�\�|��K5�\�/�B%�f�F�#�Ƽ0���Xn�I��,c<�7��T�m$�?��/�ڑ�V�*�w��NR��D%t����H#�S�J�J�� ����N>���K�,O� u�L�5�yh])C>+���{ W)��v|�c�3�٣k������L��<���p'��WdzL]!Κ���|��C�(�X�lHKz�A��.�@^͹]�6�32���`���BI�-,�ѐ�l� Ay�����]��Ǫ��m�>��f�>)����2J�%�;��(m߭�V��"y/��" �[����H����#�oo��\�Wa���n �%_k�\���;�1�N�f0hTX��X$��1��{� �I�/����"g��R5��| svM9�����:^���)\�^��m�n�f�[�>�K_�}˰9Sv��J�yX��-�w&�S*��;nm4)��Ĕ= C�u�C�ْ��i��#�4!J:6'���W��IkP4�S՘�_���-´Xx�wF�bɹ��e��7lt^a�yB����5��T5ռw����uA�DlD�4_d>�{;�����b�����s�f9W���j�������������l1 �?�ܱ��@�	���e"]�}Aw�R��;[��������b���?���u3�q�s���-�9d�~!2�鱰�Z��u����x����p}|�BA�e|n�j�p|;��ʨ�0�IW?��c�䰓��br�͎;���>f7m�0�p�w�iA��Yt���ɉ(���}'^��rY�R暇;��N쟁XG�^j�@,}κĔ�0��WG�(9?�,<����d����\��wD��	��?�K������T����\8멬c\?yA�����9\�4Ռz� }>��ZOӦS~k ���X�CG�j=�&d�W"Aɼ�P�s�[N���H`ee�G�W�j��Og���s���*����=�ɓ<2�g�G�8�S����7�8g����Z�;�DZub_�h	�6�sp��� �Cy�&G�/͘�~^[��a?֤�lӔ�U�#���tx����)LЍ9lp�Ӏ�T��D�,�V�xZ5{��Z#��%�Zq�*�d�f���ىΜN
k�5��M���|�q�'D�܇�N(,o��������BP��I,�\�E���N4fA�JBdH�	X�F�v_v�8��=��&`�Ѳ!9�A���SǎH&	n�Ă�����9\���G�l�_.ֺX����
*�6�+�e�ſ��ՙ�/M�&�V""�ϑ�����&���H}Iz��A�
kO���(�
e�5#P]g�<�H��X��7���򡈽3����-���9 �y-T
�k!���B4w���q|ܱ�O̪��0k:ټ�"6��F��	r��FG�=�JJPr?����I�������m��"�e�UQU���p��r>��1�<B�i��|E���&�F�ӪT�]�z*�t�����n�([�'�;�c��O���^u��Zj�Szg��1����t�MP*(�i�'��3~�V�π��6��s�rF����)L����~]�,��)Q�Y�-�^�Jf�-��UX��5B��D.��w��όH�=$�P��}]���v"��H3�G"?QvB�j�N���d˼��NB]~!\���y�^*z���:.耵��8��7�;\Sۃj�tO2�u��̓�J8�D>���_+���ƲS{	�T��0����"U�pi��w�طD�bpA����."��$a��}������y�D��_V�K���s-.�"W��%
�U��tPԌM���NWŁS��?�@��5q����\"�)o@�;Sd@���D.X�a)��θAk.;��?`���~Hhe��s%�׻����Q�8��o��ȣ�d�]��c�T���,��Cd���#��7�54Bt��%Aw��Ȝ��g��1V�r��%?�8sGh�X�	g
Z /Q#�}\e�t�Y��";���}��_ 8�J�]fn2`{វ�����ɓi2�Q�a���2�;Ow�ĥ�I���+������E�v���OlEg�aފ�'2Wu��E�/�ħ�������q?(��M�=��s�U�'4�F;'	%�X�+mO�tdvOm�7��Qu��_�}Hޛ�� @Of�m��դ�(��[��48-2�Z��e��%j�׭%]/�2)kX���Lg�����y����J�f���}Š�"��LE|�^xn����=�T^u �9��[OA� ����	�W�����x�����:�\(/m�}
O�$�!�ĬX�������fRjڕ�y�q�T�E&�~�X[ҳ�8:�,��I/���.�y�6�=��( �>���Ԭ�ie���<�։��y>��p�W
v�oʴ����q�pRL{�Ƣ�~@ �����ʋ,6�`B9aZ�VN~P(���_K�-7��h��J�����gn��F����qluIH�g�R�G�t9�\��k�)ю�#yP��6A��՛����"��^J��h�B�?�ɴ�t]$V�G��۪e�¡���y)��'J&��!@0]B�����(�UR.,�;{	Y���(�dx�_w�O�0��ģq�gDba$XjHi]X��wR�͎���g�H%$�~�koDWK�K��Ig'�k�m���H�Z�A����(E�D��T����C֮�'�� J����� l�Bl�4��;Q�L+lHC�����s��n]-u��ڧ1з�4�Eߡ;�wll�6rAQX��k�<�%��>/, R{��ڝ*fO=kd�2 ��K�C�D����~Ϧ�3����Z)���U|�x�ӵ�lv�6�Z�F��J�ݯ�Q�)�H�\���nvdz
��@ Z��P&�oI(.��@�E�d㣁SSy�@�	���R8��ٖ�ܛ>J��Ll��H�z�F�.�Ө��+���\%C�+��T�NF��m�t���t�*�}���6�D�H��{�^|�6q�n���^6~�b��: �s�D���{׮�Eϔ}�#4�Ӗ7H�| 	��8��e��j��L�w�������Qڪ�|�x�R �=mctZ�3�r�R�#�������g��ڪ_��M/�'�ecw�0�6g�����Sh��3!9B��y�D�h�����Cp���2�Zk�4���B"�JZ�,
*�d�$�N��v�d����9@��j������\N�.�Ǝ�k�r �%�1��wv\bC��3FBg�G�a[����]�l����l��� ��+i|4�u�ѩ�h�j�YV��"3�ɼe���dxݫ��)NvL�]�]w�/x�S㨌8��S/�'�%��8n�'y�U�!�Q��9���]o��J���?Ώ�8(��_�o�b�]Ȃ��#m�2��(u!�|�7縁�;�S�K��F-����J/>Lksc���(/f(�qFp�j�d���C����xUl��d�0X5��~_`\�?��3Aw�cl��2�L=	AA�\
{qQ����6����$>m�{�9�g��ʿ����^�Rɷn���Dz�N�R�8��-�]�Ty��}��5�����5��BЊ7.��!��[�9��[�ξ�=���-��7á���%�������S��iv��L�m&0��/]'�����׿��	��7��t���g�.CϠV����Fa�0�Wt��ډ��m���4#K�?�B�Ja����ă�g緋)]H�8����ڙ�{҅�Mʎ���@Hx��i]w�>1*ʑ_˗0��wB�}���^0i+�ϗ��e��P�C6�Ra�|np3b���N`޳/���D0�H��2�{�f�С�-Lo����qe�cx�����)h ���ff���F���|^(e�3�3�x�W��8ܡ�궯*Mg ��a��H�"�3�%��N����su�p�`��vƱ����Kc�.Li��q.F򋠉����+����#9ߐٿ�]�œ���5���뉘"�,}i
���~��JWb���,���;���l�]fn6e�����$�8�.	�"%���M�j�$�k��3��H���3������iń�L����?D͗ߖ�f}9W�B%�L�9I�U �-���#ޢd4�wT�9n�p �i�Ғ6Q�(�<;a�����T�j�z���d&��
��:ݩ��>М`�A�\	�R@�Xo��wh<�'��� ul�kM��
�İ�oV~� ���u� ߬3iBe8݊�ʧ��屉ț�ԗ@Z�V�/�5�	g�9�X�&s#	DdLS�&ܐ�/n�=��;��kI�W�5��9:��=_Չ��%Y&MT&�0�=gFS6��/ulJ�z���Y������$��ܦw̫݉�8��K�9�P�N)�o-J�h�JVsk 5[h�r䋃.�k�b�k���4�a<�$۽�q*$;(�:J2&J��"Q풞��h��+e�$����c��!���,'��&n�A��6�K+mQ�FX���3}��R�(M�N+?,ۮjG,g3Nu��ڰ�S
��~D���H��	Q�Y�z���h�/�6�n��ocԃ��� ��(?|+���"8�9�-�g,\q��H�{�ဵh1�-���!��@�yy+���C�V93..���	~ �}��dw�Szᵷ�ԯ�s�ZN��^MY��u;���}f��/X��c ��8;+1<�{*�G��)(���8?ļ� ����{��1_l���D�
�	�aˑ�D� =��m����G�P���wJ�5�U��[�#	;	ֵO�w���|�,F��jP��w1lR���2��S�;�x>�袬�� t���.R�R����/Gp;�?���7�x��fx�MI�Fo�N��CC�B!��q�#G���gX9�4�ة������ܺ[�H�w��'��u�0�~b͞�V���W�s�gk-y��.�:}��]V@��^��P�.����b����c�dܬ��ԣ0�g6N����RꀀZq�.�):��#wdP��w��b�ާ[V�	�w3x���[o�!F��:�I8�jԑߤ��A��f�錣�� q�*9�&�*Jw��lp"MM~j\Ȟh`�b��3ďT`�tz'�À���F�/�z^F_!�������N6�M�a���<��o�S/oE��;}�;o[�Z����i1�a�)J,4ʏ�Js|�q�/Z�� ~^+�t;�����tW������O��QMf+�-C�	�-X��R&���]�,d�ʌ`������_gnݐ�x�Dę�f/4&�Q��r�C�3�Z�?�NT��`s�Q�.���":��1ڠ��g|�����S��W�|R�@8P��-������������*3W����L��(�M11Żq�w`�.�P���k!�3ܚaQ���G@�&���v���:aH�*31z��^N5[d4��^|��t�).������8��v��Cg%^R�"�S9��	ϳ��Zq�UBe����p��W"�kn\��X����#4��hi>�$+��D�
�2̀�?�?�^�:1�)�@�)=��WۜRҚDk092��}���3�xd M��qU�,1
�uޕ��x���c+.�px�ޓ*�2�T��������h����an#�Ȥ+8]���Ŋ�ufC����A�]r���B1񌬍}s�KV���D�$`rR1o� �Z�����Q󕬻u����r�!�	 <��@���'Б�,~�D�
] ����t�gHn���3��J�ke�"�e!с�z��ѴG���SrP�\;�eݥ�,��q�~ �@���;�����%�{>���)/+-(�=�����'�ܷ� �}���[�/�lT�3u����Y���������ކi< �>��Y��n0B� ����/kM.�.X�h�z���	'��:�>�D;�#H:��
$����T���ˎ��}�1�1��]
��tch��҆[�/^�3���� ��|�ixQݔ(l�G3?�><�Gr��2��
�7���M���/iv���W��>�Zr=��cs�i�� �ʵ�������U� �������T�U-��(nq%��)���MoD{���˹P�S�az�K*�K�Q���PACU��Lg�Ȉ�5�DCE�=�(��?����B��E�2{��b�9�7�2�����5�=����}���Թ��V9��^Q�$�c���'��%���6G��T<��|�pL���)#�L��
ϯ6@2G[�xvg|�PB��0��IM�$�3�ٲۄ�]�tE { R�������A�U�O�d ��t ~ZM}�f e���F��
�.��$���=���N���>��Nh�D9�j�drg���i5��Q!��E�	�*k�Lx��1G��趟�!��H���>&�*�� ��c/�9 ��n�~��^�^�ψqM*�OE���
z��&�
�*�b�)�_>�K�j��qy��n�"�����N
�|mD�C7�)�Ȱ�ZB�ş�a%Ϟ�{���	!:��������#&^]CA�)R>��F3��� B�?;p��Oޢ��m�C��&]^6��ɯ^��Փ��'�7���`�:����{���A�R�W���������,��
������$�o|�/m���	�������,��T�8UX1���~�;`��#�#�T/r[����G�g��0(�ܪ�!ka����v&S/I�V� j|U� @D�fG�t��OpR�ѧ9���Ȱ����\"�uc�6��a�C8���z1�7��#%�k��Xnz"�1���^�f�7X�׍F�'�?�T�-��RoC�S�E�"�:�j�!t�'7�Y�p@~�`�2q �N0��P�ʊL����s��/0�.���I��'��֕�tE���E}ȋJ�'5S�"�n�B�����"੶P�o�	*#�@z�Ǥ�Ye}��c��!ZiFK{ґ1�FA{;\2�sy���I2K���B�+�ڗ�E^!���}]�"4��b
�E �Y{�ē�u>�b����aE���&f����	����� ��u�z��a�����c���j�j'g�eS't�7���\��=��V�^X "L�σܢ�S#\S�cd@M_��s�����9���, �sl۰,>(hF�����1y/��ɜU�?����bÉ�����ė�?j�j����TF����uR�E�<��-sHYg�����>侒Ϋ ˝i|��.��L�[]��Xᴴ���K,�����!(�v�e��&� <^F��q�ϱU���f�����<�G'g�5�J!��P?"�J��հ͝0>JUY��yo>߼��s��*���9|q0y��9��d|��M3ٷR��>�(S�#7�޺'��������^�˹}�+5�|���6��i�0���[A�,ls���Γ*{�;O5�"��=鱛�U��/��5�J��f�I?)�{�8���9� ��#K6|��� WT/��`m)2�E/;�x����^E����eÿ���a��V�S����B���:��i��,]��Ʒ������Ƹz�s�"K�K��,~����O9E�W��&����<��	cL:���zBB-��Y������ݹ��y��N��wI� B|�j�s!T���W���(F�&w�O^�k���-�%��i�mꜴ��do8��k|l|�I9|���J����wkL�Ά�'�u�X�0ͺ�jA�%w��?��U�#6(�UQ�aH	2��f̚��6�6�=&8��{��_��(F<�Gh�$�����P�P���p����Rf1�L�Ҵ�a,���Eٙ�\-�}���u�Zk��rT�Ko؍}s�dk�91��[p��)��q�˰>����&�X�3��z35��&�c���D+�{���6{��DD��gDIAB�Y�J�(��m����"�A�g��J5I��O�-[��A��H�?7u"�xI[�����m�8�2�3	?a���C�b�v�n���kg��:/`YO[���~N����h�D�D)�'p2�&�)��~�U����.���"7N=�7�XN���[�;��w���~~��*��:Yr瘬����sW���G)h�ދ"�,m���mo'.Z\]��	]Ek=Ip���C��.Eꆖn��Y/=v!��Yn[~�x��n�F��(k��;�!?S�����T.���/X�gk %G�svTVo59U��)�M��˵)�NM�}Һ9����w�`Z�c�_���mK��"��7��xDu��Gd~%��s�z�����Ej�d��s�j�,�#�-X�dd�ds����������|���+*R��/�FH��R�F�^/ٟ޿���y³���'Њ"8�5:�FwC�F��տ�ݟ����9�{�������O+ϳ5��2��!��ʟ9��F������@@�3�+X׾I������?B���yG�ML�2m3y�Q�2'!�u����9o�GS-K�S]�:]"�`�V�T�uH�I�V�	��s�cMj>B�HH@���@�e�#c����Р=ł#�1��a�j�>ѣ5��SM��Z�ĉ�!�B`�$Y̲`K��i���b���;���[Ʒ�ڲabӓ|�x#� ��L��>�P�K�0��M��!�?ݙ�H(�a��rh�Y��G�LG(��)h�#�M������K6���_4]/8��'���G�H��fP8�J�s�Y)�������M<��X�M~ ��|�z"��ؽ�`VjX�3�Lm���;x�z�B�2��� t|o��gR�����y��b� ��®�(���+��弋��{���
��1�19����Бg��p�bP`~}@I�p���S��D`�2TzV���7p�_7�S��-|Z����7'y���h�|_�
J������@�4o/3�9L��/���{�s >3��6<I��p�8Q����Rp*��1X_Ĩ-/�ﵠ ��;�o�ί����d�{��*�¯�|����>g@�k?������'M��j([ˢ��Wxf�%x��{�`qd-Y���ۂ�xtZ�S���d��j���v\���`Ư"���M�;M�� *}����Ls�g�T��!p㰬�}|QM0�F�7��ӈ��"ɛ���-�3E|+6Ѱ� ��u�,A$����O�,"��g�w�Yz�Jf���s0��E�H�击��W?�,mЊʃ�����(>���q�2��後�A,UXj���P(E�*e��K��
�����k�s@w��!;7�S�X������x�Ѷ�1�V��%8��%{�ʈ��)n �M�������>`Q���s��F��/ ��=3Ԇ��:}�*����\���\��^~��7��Cһ�^��L,�����Tv^}�/f��?�sӗ�-�U�DZ)��i��=@
KC]w�i��1�$�J����D�ol�����#�S�淍'������mc�FS�:�,�A�	J(}�XDj��ۘ��bV@���ҷ
c�(J<����0�!�}�IxSh�p��N٩�S%��ڼ�*�N�VCCߓ��u�4��7�B�Z6Gڶ���0ϖ�}Ȫ=�q���'���O���Ҝ�M̸(Y��Yx�������Y�yR��׳ږ��b�dA��4�ʀd�����]�e�ͨ���a��l�����:�fb�I^SYn9����֫���ګ[�:]��Q�cCr���X�R�孻��������D>���?H�*[��1|�Ч�za�2Eyb��w���ou��D������V����/ph�X�\sX�1LW�����Ax����BV/���m��;�(�'c���%N�d?0՝l��HdD|�8RMM�k�R��m� ��T�a{��1P]������Z�\7@�w+۸7Z�yJPeqW/�1�7���.�Vgp���Y-$э%GݮȀ�@��\�87t[�=|�R}MP&'gK�̂Qv/��o�ykIc�\7-�I*�?w]�͏�W�c��g�ȍ�f_8����#��,��-`"E����X<_������4������q\��wgB�k�k�99oxlk%�9��3�
#$��<����՜��3�{���ɢ����u����K�iC�s]��W���0/�џY��0��|F�f(E����JK�$t����ߵK4.�ÓEzs׺O�c��MM�������1�Pb�LT�et�9wo�s�f�m=�^=��0z��N��-� ^�^�Z���ޗR�R�@����R|cg���i۷Yrd1gft\i���U �9�1$�	�p'G��{�$b;[,(m*���W�umՈd8��aV��Q���s��w#w6Ȑ"nY���r� �{�l�p���g�U����8��5~µ4҉�y�f.#���Fʱ%>�Z6z�(PJs���K��B0qj�~L�2~���$Z�B��%��rY�e�j��XC��z��b��Q?�|�	5�(���:J��b�ͼ"Tz�X/�_oJ'n��� Z
�@�/���%eە��fg�
���6�,[%�7頉p����X�o?����尭�ȜA5�:�#o�����
!MA�llٚx�s���������!#��K�5^e�:��ӱI�SG�Փ�<������ߒM���nYʸ�k��L�^F�١/��Ua9Ql5������!��e� �BV�_$�;�j��k�?��L���N1��p<���*
ʶ�z�E����V>N-vM~�@R\���V�[Q}ZDޛow�&�8{�����ي~X�H:a�w�{�3P/� ���y��E�w�Y��;b�b�*i��t�_64;��e��`AQD��1����+�����'��@�U��@�Z��j��JX�g�G���t"�D<���R�60���6LO�M(׉����;ϊSEcF�vQ���C��Q�%4�V�bZ�.�������$�a��E�;�+Q|I��z�vw<lꃲ��2=��)t�2u�x~Rea+d·��JM��]�����'��xp�����:�p=!��J m��*���Rb�-c��5����S��rөk%�j�#nV��2Ed-D@��ckg� �#B���e#�Y�Gg6�BP���"�	���a�8)+���
&Q�����rw �W[����Ց��ځf�LƁ0+�(� ѯY�}R���	�	�;�w��8<^`��8;(��By�Q���59�J9BM�Fv~h_�j��.F�{��[-ښ���C����+� ��	V�_�[Ǥ0GR�(��.t��,=�I�C|I���	Ծ�$b�M�>7C��9R����Ω3���SU[{����p�k��ve_Iw�����r�h� �)E�hlԝ+���a�풦]!�������e�9\I]~&Co:ԧ�a��)%�G�������;��@��>�w�n�S��]�I^�x\�Ȃ~ ��ҷT����� 8���� ���;����\�<��=�k����9U6�$�ٗ'�K��y�	V`Љa�^B��e�#h��<�*H����T��Y�}�l�]��oA{]A0���Gn�Qjo�d~��o���D��,o;4��uԭy�|K�)��D�u��(��a���߾�.Dm��T�A��B��Pw��U���)W��!�U����/�ĺ��	�����:�~��D���}Iq�x23�z�V_�����MJ\A0c�ę)�OF��e�s��t�k3ga��v���1�C��4�%�9;ζ��L0x�+���r�&Z�ۍw"[���m3��B�{@/>X:Ҫ�tꦃ�tދ[�|���R1�=E��%����Y��
*.���#��b��nBʞ�@��������J����!{�����nf�0���VhH�5����3j�%t�f_�A�A9Hq:�̝r'{�ۓF�Ak��C��������(X�vG�M��,)����8J~j�	d<��X���ΤH�����	Hg�f�`C�X�B��>�8T�$�L��jx�f�h�`�w�vZa��I`�	O�,	o�@A��e	5P�>��Y������N</���Y1������9 ��B��<�Ig^�k�Y����+2_����4�R=��i=�<q�)�"R@ڈ����J��|C���p�#���FM{�J:!}b��G�U�P��Eh�Y�@����ϸA}\�u9�r���EA�Gx�&�3��`��*�f��=(���.��+>~��ب��vO�P�ǖ���%���W��a���"�55�eb� 1���d�q83+�S�4:U���_$Fu�Ua�PA10���:il3KB��W��aB/�#��Z��ݭ���B7�DX� �I��!n��[��-eg��X"4R�H`��g�]���͊bn�06��y0L8l0!�������Rb�!�爸�ޒ2q��}���r2}iJ�Q��r���R���PG�.�^�j��RF�m���7��zQ���S_�^�F<�+ˡ�g;b��g�aL�em�eQ�,�3� �&�qf�Ŕ�īā]tm���Y𙐣W��|9��iz���ɷ�v�njK:it�WX��PX��V�a{��>RU�5YaWK����,�']�'p*-=��4ȳ���������w� �P���W�I$D�N���B�M�YU邈9��<i+�C.�yg�km%\��S�L�B�����ԟb�1��O���r�y�������9�劮����I��wh��f��Y`�80�2q�C��;�ap_��PS��v�c���@��81�hO$��\���d��)+�;�%a2��)��q2Ǡ�s�\4��2�3X���]�<�%�e�P��G	�")�c��y��N]MY>��Qpkc��Z#��P���έB��kG���ڵ�o�����R�G�^>��S�+߇'�,b������OD�<Wd$ts�w�7y�JS�r��U1����\-��ЛugOpA�H�.9�^�9w��rA�5K�o>�HF��@#����}�K�5�Mꀭ�@��{CԵ�ׂ��������n*�$�]lq�:��U]�-����
b�d�S�e"�T���Pd, s���1qZ-����Q�K�eS�����r���s�=
���cMRfGK�Ԏ�|�b��2�u���e�/:�f����+�j�p�W�	�k��î����NT�`��P�����}8���.��&��Z�ȊS�L�L ����Q���Ee�D���jv���۵Ѣ�z
(VyW�D�h��US��[�\��&d���<��^�5ȭL�ћ�[yqԶo�I���KG/y��)8�������T�^Q�Q�[�9-���@�q��Z���������g=����&�Efov� T�M�����g��BuǄ�1�l�.B ꚣ��]rc�\o	N�}�&��2>��"�@�s�೴������.���.��Ln� �;���sщB%��p_�����US�-��< � �!F*>:�������lA��Hf?�����c����*�p�}�`�yuH��d���:�����o�<�ҵ G�#�?������j�Ű��
b�b���fP���� �����Mxrޯ4ĥ�.`��(n��:�C�'�b8��N[v��a�ݶ�T�,��U܇*]���b� ������ԛ@�bI���e�602�ϻG7�h����@�)���+�V�	챿U����U�v�5on΍-/�B�&�Z��t�+�uyO�>H���WSvkb)��!ԡ=���O�@�ö��Шs�p��U�v-�	��ۘ���@'�C�3&�`�������t���[5O̵��Εc��k|!�37o�e?��5S�$���0�0��d�j��4�؇wL�I��yj�E�z�\|���v-{��F� ��4U��/���~� �)�\�Y�f��#�7Ը�����$<ʟrh"�|z����"|=*۴󶄩�irK).m"��0ʖ�+s�|�&(��h�g�L�FX��hl�&�,����G[��^ ��ӡ�'Ҟfë84ԍ��}s�)�����g �?�>6v3�X�Z��Y��P}%���O������ov�I���ŉa:��<����1&^��b
�D�6��<�$P���*�4�����Fk�Bî��,�:+.�#彾����K�XW^�o$49琩�Q�o���J��t��m�!��~�>�.������w��y�hU-��3I.v�&����X(�DJ�&ʸ1J�f( �s��(�C�B��m�n�¨�T�G�t4�L�7bة�.�nH�Y�ji0�=�F�zYd*�jT�>)�A���[�x� V�[�d��L���-�w��R1i%��Y��:\�������u�y���,tT��f���HM����q���Ρ���i����b0����S��#[�c~�� ,�%��vS�3��_&p��^f`i��k�o��w��{��'�<��*��b���,k�)zq�_l��\���Xlo;�ׅ�J&d{���F%aS��@&��*�p�/�$������]�|����9d��� �|FZ_�#�ǅ�g~���X��v+�[�>S3�9��`Y�����'�]K(��޳բ���C��m���dԼi��N���2�_�>�OL� ���p5�a� ����S��:����VT��
��8���eh7�'>4
ȫ��C珌i3�]L�� [v�KuY���s�W52�6�?*��z���Y��]��w�|齀���Jf띾�:�<���������#�"�UF�P��fyRq�
h|Sb�F4�#}I|I��cQ;��_�rdy��d����/�l�沸s�
T�ʉҧ^R�P���YڦOS+D�l35s�D�׎�8gx5A`�iH@.�WĵBT��`]���Un�;�V�;�Ǜ��>�G�RNp��X`�+�=�Z�?�Ft�?3��/�������yP�4��	���Νs|7�}���X���6��h�����IN!���)c��N�-92]�@T-[
n�^�n`K�T/ȴ-o�%-/=��&�E�b��rb�X�y�36=�i���4�H�����K~��S�8L��$�ö�!:
p�0d�"���~Iܶ���f�p�(�Q���E�:}_۶-�m�
Yr4)͓�}�!��)� �sP�U���PƲ���9J��m���M��={��#�2�[�Sr�ql�4�L�Y�^��O�<w���F4ґd�Ǝo��=�k�8n{�+�Oqc� ��o^��m�OC/��~Xv�5C���^� Eȉ�4��&��8�l�7���"���|�cR0kcP_���!�(,c6�M(�BELIao�|�����d�č4+84���d$%��Q1�ik<�2��\��L�TS�	Bv�\��`*j�[67ە�t������ˊ�[9�"�Q�V�@�����1��(��翳�h�Ye�	�Rr��vkѸ�&�0��:���l0�#|ksP�G�N"�D��]�Q�٩ s����lx�-]�� �a�nZe�<�?j8͢��AǇ��Ql�ѣ�p�2��];V����G�Yw7��m�$�2p�>�_|�w�ZB���>׃�!c��YbQ���~����
$S��̸��d�P5�ͦrIQ�1�{2��{�#�Y#�����D=�������}��d�Z��j_HfM	%�>��O��d��(DM���E�S��.D
sĚ&_�6=��I�e��z��f?����{�SnѮmnc�{���;o�cf@B�9�KQ�㡴p&�2���w�03W���F��4�o`���;c��k��I�u��o�F�ҕu-�Ι4�6އ�����5�Ɖ�00z�ͣ� |�Y�kBUw������i��T~��'�R*�����>�fZ���3�֞����=8K����"Y '�,e��vx�e ����)\<N��������s�|�I��vIp�L�x�D7�_��OJ^'�4=��E���5!n,bA��\�Q�'����b��~(&� �E��]��!A���
Y�Zшyw)�n���6$ٚm�c�!�>q�])1�h��<�S�:b�\'�Ad��� Y^2�?���G��_��]R�'���{qE��������.܈�A��6?�C�OP�� ȭ	���M��KZ^��y� �Q&ˎ�<���?G�nDb�c1x75�t���%�W7p�I���'q�L��2$����y5�k#��r��h5�a�Q�t��W����>��0��-_i��,5Z!ѡ<�B~뾆2%�(�z�eEK���D�/U���U������3��۔�+�� �)�8��@������^J�& !�U\,� :ZOD����P	�.��2��a7�r�MZ[�1�)�E���̿s!'B��'�u��=�X�����v\-C%g���jQ�?j�� =LWl����de�FZc�~�E�����>]'�lG����>�ː5$�<��HA�W���I�tt�V���vERf���Ґ�tj�{8p�/��8�ţ�UjJ��)d�Ur+�Y�$�,�������#夒0(^�u�i���;�� �y��j㴪#G�Ɣ�a�e�LI8�zD��Z��i�6S����gu��>��>�.��D+�c��q�����۵���H:{_�F���W�^�ߎ|��K���w�2� ��'|5����4d4�^-�1��
k-��H]�C��U�������lŏ�5&����bz��:A�^�I���F/)`���n ��
��9}�_`A0��\׶����3L�<���dj�B<�tE7V�LKLk����ō]4�ex��J;�0�D�fŮjTc]�<�	jY-,��.�K��T��C�V�SR�p�#�Rܑ���qFC�@4�Lҁ��]�ʓ��xz�C�E�#�W_ ��C�R	�Q�u3{����(6�$�e��\���`���?�quq�~���b�%!{)���C?s���|�Ӫ#������C�C�fe]W@��:2�{�%�M��4�L�Aj%�2����ɓ�4u�Zv��ѕ��nfa����CK�4�Y�Gb�q��r�J��h8'����wZ ���9��?Jn��e�Y.�J��' �k�~��O>}����-��]��q�F:�`7�D�E�f{�f� ��3փ R=�7?g/���dTf�^5��*�9�"f껬MCS��w�d�^H�{������!L,ֆ
���U����*1��?�����"E���a/Ta��Ց�3�X�:�"�a9Ԍi���y��ӛ��"��?3�qF7�r�9�q`�;ť�4��)箕XN��[:��ĩ�\���=P�=s�%֯��#]��dQ1�-:i�����l��	����Fu�����T�ݡ��Mq�5v�'�˼#�3㏭����<F��N��L ���䕃�K���h���_���qf�L�~�u��(�f["f��|.y�1R>S�����.�2��$��)�8G���%��_���)]�y͒*�"�Xj�iȽ J��Y/�9�R/����TbF�����WBlDWMt]sV!Uc;5�lh9��OR���|����^=�h�J��RL��[��_���,����rŉ��,����Ҳ�-�tK�j�����t��7�=7z���$P�1&_�����o��u�
�?Q�J��R���Eaо��e����������o��8�n\j�}��
	���il��)�r�Q5[����\f(+�!��qV&��w�:�\K��cr-�Q<��������믘�	�<�3� �\�N��'�d�J^)�P�k��1�G�E����WT9ԑP�ZS �Z}��Ŗ�sr�����u&l�ø���JZ�K3S�}�������&��Ր&�}Qe���]�#��|J�˕Λ�{�;E�&�0䟜�O8�T4؟
��E�d�����>8W5��B��ѣf�|��U�YNf�w�?M��9m�2L�L	�mPr.|��cR�a���dޚei�}s���-�5�޺��Pf����2��)�V���/D{�n�޷$��ܹ���w��[�{����$0,��f΋"1���H��6E�$�b�Y�>��ò������I��Ϊ,�iI�b���4;�ҵۘ\ey�=�_p'��K��vHȕ��qDF��ӫ�R�TH�����#��s"�j�*�N�t�%^9�H�L�ui�H�|�3dx�$}�bz$A"�{P\��UK��K�a���U�����
Oa�yݒ�<�#Y������7�R����[��P��/f<q����馆e�+z'Po���<�|f8k����D�	���-l�e��'GP�@�Ӊ��/W�R��5��m�"���K��"��s0��
 A.=P�Q���X�qB��*��GR0̕bLR�
�f		�g���d�:��Ӫ,��p��rf,�xzb��E�9��S3��={�a���fNK m�b���b����w8K0���=�W��Rc޷/���H�4����b?a`�<��ЉۓP?֏����A���l�-��{AQ�9nQ
>���Yd�۪I�d�?��(�4�0���M��LrZq��A�� ����NL`�hD�O CI�XZު�8�)>�⊎����]�@�k�WqB(P�5:��O(�p�Gur�>��R$��;��W?1�4�(�C���/0� ������m�8� J��;M�=�P�r��T�6��x�<�TVsl��1�.�g��?i:�C�z�x҉]�T"8ba�I�X ����XBq���r��g�!����$��"
'�(磅���k�c1�jcI�\EQj����ė
��:�+M���tp�ϐ�~��fr�Bɹ��t[�(H��,`��,hå��Yԇ��3
�&�2�a%��}�@b0zIך�`RҝcYn�y5�i�X!�"�l#������m(�M�����k�D�S�lvNVP��q�0�6x��g�\�n,��?G�[2SO�֤G1;�6I\���]��_k1�)�Ȩ�
�!u�S�T�v��+G�F1T��jE�ؘ��U�oj���o���Y8��
4���t[*X��a���Ҽ�$Sl�D���l3 ��)�}	�vH}l���敏�l�[��v��2XU<2V`�l'�w�Jo��.�)���3������I�	�!s8&.�g�\D������:�J��t�{�`�w$|eA�E�q��$8�{1H�eTK!��"��i��U�'���.�&�_�h��+M�D>�.�j�
8���L�4��@x��h/�M�z���ii��v�&��A+V�V3׏�%�k�9g�Fu6������z����׳��剞hq�����Q�"���$�h�_zL�����o����BE;�([�j��3���	�E�ğ��`��z��^ิ�����r&���뀈
� �ϙ!Z�i��z8��7�m����	 ����
V�fPU%�JwhҺ�z�c����_���I�	"�0C:��)x�R�$o����CX܉t_ V1�Ө2�6�W�E��4�y �����a�r��S�K�]}G;�{�C~��a��?�	�|�D��x�Tm��rr�2��Jd����;�P�q�k�z�S�D� ���b��j1�#�B��O��UPRȅ@���8�^������8| ���	��Tz��)�T��-�~��7mC�Â���o٩о �gR&�[�e@��e@�+��!�}^��~��d����t0�X��P@7k��^�e�,�J2��D��F��zwU���j�L�'q����h�;b�S���j���Hn8�Y�ic��,��c��6�y��I�]4�|�V5`�t۔R��PjVv�X���*�v;9���n~*�܅C��o��iذ�Lb۠qhd��p͈n��я���5٥)i�R��I.��x���A'q�gK��U2aa�&ߩ/����֯T�y&`h���FVZ`e��߈?%,��1�vN�y
#�sg`3�@����X��C6�|�g]������r*gGTG�s�7O��|��p�����0B=���5�1]���AM�R¡6���8��S	(Y��Z�}��tx�!�[Bn�&���`�	���&b�6�y���L=���S�� �G̈́ۗ�)V��阱�z�(�l9�۷��F���F�:��@:��V��Pn;��(@��`N�7Qh��*l �W��An[�CI�*FUcx-Z.�N�/�<�����t��R,୿��h��-����D:�4�K� ��_e$�+�}c��0(�SW��G�H��U�ꟽv�����s �����U�̗��m"a	���]���U�r��s�)�#'��G�:�O鵏�K�������yD�a�k�}ҐE@R |,D�K�֒���������� ��T�h'M���I�Eeg06��7�(ms�Q����X�&Ŵ<���ܓ�Qzq;��<i��/�p���w��` N����VM�_0�G�jN7c7�yKGm�d3w�K�O��� �:Ib/��vO���)bUk�{�i9�����~��I<,���"G�J��֯>Y�5�1�jѶ�F�|�faf�����2I �/^���q���>7-�&� �	�X%���`��>�yHQ���F�+�G������?�NAc 4�{�D^ZFJ��,��]�0�".o�x�i�O\����۾rG&�>nX΍��K�l�o� k�(�~� O7�_x)�E�X��,�I֊W�Q: W$w� �����O0�O��n�>�Uo��p��2UX����l�u�:�ȰCB�,��7�3aۻqSAl2F�#��4w���b�I4�}M�?԰@.�?��!�A�tʕc�; e�Ǫ85�^��A�D�q)v����Bs���Z�?Xe�/76�ɣ�"� WB
�=񗾙��|�Y̞l:|h欦'���*��$� o3��*���i�� \�����S"�_a�[�Pk��o�/�����g睳�u������R�D6�~x���}��Ӣ�1MOַ�	([~0Iz�>� &e��E�p�g��ƃ��W�"b�1��O��V���B�zJ��RsW0��~�i�5a��i([��Bn1�9'L�zd�:G���������5�5%��HRl�ϓ��N��ri��"�q��Dڋ��T�:����b�ԛ�p��kU���Kw��('U�j?�@��L%�:|�xRj�+�K������v7	I)}[��^�x�ID��Z��ⶣI�S���Zu�]� �p�.i�]��Mx
�
)� ���fC���]�+U${�T
�.y��7#���k�Z����d����H��J\0���O�2���Hk�d^56�].��u�n;�~i-�(c4�e���.U���c?0j�CD�/��6,���L�`9BD����@����>�,l���1�D�\+�VC��s:�H��!`�[�)U���R�d< 鼂xcq��u���@���L�$�*YO��K�(_���vy��lU1���Ψ>�՜s�ۯwxrQ&�&� Z��"����YhY�B��~�[4���q�m���.sCU[�5���h���	�]=,5-A5�<&U	<��J�u����#<�)m'���wCƄ�=�8�.����?6ՙ;�9
���i�n5Y� ��C~U��f�Q^tt_y��`'v�]̩��&8�H���Vْ�������,g�#�vLlN!R_Q	�$%�0l���:ƛ�J����'��0�}�zF)�t٤����U�K�4p�2����=h���F�R��哷3�3d'R��IrMh�D�4_�_����.
��c�������d��G�v���X3��X��G!vU�߇3:$�K�v�xٛv��,���"��=�..m$k$B�!��R�p�%;�{�L�:�1�6��j��>d3����X�f�M=t����z&QI%����3{x.S��e|a�]��U�JJ41Bt�����U/6/��PܛH;�2�;��窥2ib�!?1��}����9-?�]�ɫE���9��>��M����R!F͝�\E��Tx�ܫ\N��r�7c]�x�������<Y�U�`��7��˭ʸy����x�7ٍ����w���)׷��$|VOت��%�\����_m!s�(
zt5�F\��3�H�O6x�.~qҜ%��K�+g�� ��=u紝�Q���=3-r5�*�0xd"�%xc�&�1�����w�r��B�}F��:Zp���n�X���N/��J,�U��%��޷g��
^E���-���]Wm�	?"�S6g���%o
A�[����$~zM�H��B�S�B�{�S �8X0�u�:�ҡ�d�Π�&4���Fx�6�iDv����s�����U�o\�h#�c�1a��#�&�6�q�������S3�U�(��+�d
OC_�g�0��e��C����U��h$|�=�GfZ�#_��+]��%e�+%�wRﵑu���kD �zP@�|>gܮc���N�Ҙ�`�tDSN]�� �ٰ�㣢V��ߪz$��� |�X�����xin��![l��"U+tꋥ;F�aƘ�F9�b��v�W���Wn ��L�m�u6���2UG����04���iCzV��@YӴ9YP���]���fi��&��W�n�͓�f"
��C"t��!qFv�]#�m�RF���!����­ö3*wM ��v������L \q������rW�p�@8]�~���T�X�:��Q�ה�R��A�z��8_�=�pV9~�b�2D��b��l���[�T��h�\b��̺-��O�����NW�۪o&��֦�� T]�.�|2 i����]�G\z0�}T���u�F�X�T<��Rz�g�ST==�;�^{��I�@@E��c��TR4�Մ��(��D?�?0Cfk%�n:�j�/�\�Kأ�Y��~��@]��5dIB���n.
��BP4��D��5������p���J62�:YG/!'7����&�ǹo�)�)u�
�̆Oxql�f���$�Ａc*��w�!�_�.�uZ��-Tˇ�������eqɩ��� ��D�t
���;NS����C�:������)	J(R��U����E[#F�L��� �"o�U��%��;�≋R���pnѐ����}�ε�-s7ྎ��rŹ��Ɂ�nQ4|��pM���W�M��h��E�@L);��b��"3(��%��m0j,v�+;S����g�Z�٧ ,�0�^J:���B�En�-1K�sh4�Qݔ�V��Z��:�l����6�Ѳ���k��K��cW<Җ>iK������ϖ������l_~�Ӑ5jyb-�+X�5��͕V!	�MD��'sS����~~�.��-�K�[�x�G� �0*@�߅���]?B�L��1��'Oc�3����^N��Gk�L��k���?;�B�H��p�B��_�����Ow�j�I�&s��R��堂
$?6S������u�KG���	���{:Z Az)��zp����L�~����� |��n'����2���rEܛs{Pȶ��&1��������C�^Tω�!ۮ��5x���Z\i5��Ś��N%���1��zQ̶Q����<�뾺��ۤA� ь�G������H_��N�p�N,o¦�cr��:�a|��$!�������pЯz�
�=��d�:`�W�X����}�,Qn!�Z?2~��[0�r���?�f��嗀��_*EP��!G���n�-+����GP�k�Y�c9N���
>�'��Uo^�ḖI�4�Gw�B� �t��g��H��K+g6,�E�ߪ��f���w髝���9�)pV�\;5)J=:��*#�G�%��L���+L��#lr/�ۍ�HU���:eg�����I�,P��'@�@�����v0S�}-#^����)F��Hԑ\!��Ө5��h�=�$����|�����t�u�!!���*��^$W�@YE9�N��f4��L����dg���NwM��!��0�E�{��ԧ$�щ���ӎ2��__�û��l�����k.W�a@�Gh ź�J���OtWR������Ӻ��< �G�9~���7)���'�?M��e��}_�B	���|�ڂuE���C���Rl�8��s�t�H�5�OV���m��L���Fh�Sjh��n>���ſ���n�0���2+�!�tr�u�]�܉�4(�X�X5�����'!@;ho��5@���lP��c������A%1�b9�R]��Ͱ��b o.sJGכ��E<�n.7��<����9�P즊!ݐf��<��e�jgXq��T4���A��:�n#E��j>�Wy�$4�z�4�S��9=n�W��*%
�emM�r-�8��ڷ4��;?=��1��^��� �I!���jϺ����y��+�6(��"Vqa"i �~%�e�xq&]���͈����+�Z���TS�و�kq����ۢH�d>A����΅�u��GV�ڠ:^�ED��܋f�����&��Gd}=�vT!SeQ4)���{]Ѷ>Y��bS��,�
Ac�ec�γ�-(�������A��b�n�z���7��#f��xƄ@����_��i"����⼼q�q�s�=��ok�rb-I���V�O�r�����t�44U��ﮓ�e�W��6�4_寭\U��ZI@.�2���rRԢ�y�ʋe��Ĳe���?!c(;����i/�i��h�4�(E|>��l��?R�c,�w-���4.I�8��!xcg��to��в!���1�x�C�g�)�Fn�g?9�]��.�'4���у�E�e�8��
����$�x��6��?�iY^i?�x>�7�
��I�/����,��|:�*���z%L6FW���	�y�6X���p�4���j�%h| ^N:
%�:WQ��3��sF\�[LE ��~8���N���4��	^���n��h7)��L��b�G�Ï�IܸLQ�V����f�,m�,�;TJ=?��>2��i�(4�M�Fۨ�U.7����=f�+mȐI窫�30?'n��ca���&��� &(��xx�D@%���V��]��c��5@�C��Pt���@�ϑr��8y=��m�]o�ț��:�X\m@Ջ.+��U�U$���S!�
5o�"�4j 7�o#������%T�A���s�kH�6c�HJgG�����/<�d{KM](�x�a�PA���ht�_Q:���%\�e��/�J�Ǉ��)���`�5���q}S� b��P��F!_�Y���䰐�oܻԀy�B٘*�� ��?�E�v�f+��46��q�����N�r���= �����<[ifOc��;��{g�d]�{Z5!(���)�-C�$U|^�aNǳ��
�.�kܚ������4;�o�P1-�@2�Q��E2��M�<��\aj�&_b@r���w<����EL�J�%đ	�y��ml;>,n7��.�W�Ɵ��kL*8�;.�՞��=X��2��|��7�⪢�(zx[0��3�3�o�&h�S��'$�@F*,T�/ a��o�gC'��7C�)0T�T�k��q!:�i	_I]�?W�����Hk��£%!w2��g
1�J�5�w�nU�bt�""h!�����nh��(���ƃ�g>$�H�I�h�Xd���a#�-y⥖����/5��;����w�Da�u�����������1�B
Y]16@|�e\�O�d���6����N_�T�1��W�5��fڲV�38
x�t}��+�����ӆ�������u&���ңD����Q��9���l��b�8�:t���-�ck�S*�z�+]�mZ'�u���7���<Ă�	�2�H���ՏE�����Wh�%�N�|��O����ENL{��� ������.�͕K8��<�4�����zi��\߃�f����Ց�Qn'_'w��u��Nn+��Z�a���9kd����u�uܤq1%&�EI��?j�:cP�@��YۈUSДG��\����V,��L5�م���yp�)���~��R���c&�G��(KI�m'�k�gέ�c��{
�(!�W�b/c� Z�� ��Qa��A�C�[{����B+gj�%���)`Y�b��2��#�JN2� %��G�~���M$#���/��VbV�FS�V���Q������	0�U?��L��u�b��;4B���'���j|?���3xTVæ��1����u����?�1��a�����ƽ�X����!"y)K!�M).~C�T9�Z�9��%{�?�K)pp>�ӑ*��ѹ�1�V�tDU�3[hY�1�2���E �L~�)�Cs���������`�u����(ߺ�<�[���O�	Ͻ�kl�&��8��k��!��n#S_��k4���e���!#I��y���fܠt��j|*�Y��6�ǫ	;�,�%�,��g`
���h�i�8����}絓���6G9=�O���ߺ�)�����1��7���N���1�v4�D	��`���S��X�^��|p{�T��ů"R�ڏЄ�����%�+��	���6&"���0�[/�Ya=�.0�y�8lo�b���D7��@�g���VrB�/+__<>,���"�����|dK MF�,F"��ˀ_`�_�� ��+�gJo�/��\i�����O}�^����>}e�.:г��ع�7�(\�n�׈� ����:�m�������d@��i��0�hY���Łܧ��kz�	�N�qM��i�^If���MLMD):��	Ɗ'ڕc��˄�3,\z?>A���-%��*60�����*�)�,���˅eG���a	���EdBY���hz=7�J@!\,��O�1�x=�2m��UD��uw���Uf��ynnE����B&���=����jőxB�t|
�L�d��$����31ɖ�l�����a��~ck�П�~�PBd#���X}�R�?b�GA���2"�dh:ޭS��M���RX!�` H��9�U�ڧ��(m1��?K������Z�Y�J:��"[u��G��H���ý�h���&���`%��/�>��\��8���C�����t]��pt�򊆌{|%�J��ș=�jӵ�B���I��V��K����	s���_��3��d%L�7�oP�����T,���53$ �Ѭ�z�'QhI�S�V��nEp��fm��o��eւ�B�����B��]�2[|P㞔	j��s$Bk���f#U�������e^���P̳WS�>�^��ض��8(%��6���[�� N�&�\�{�5�U��Mp\F�5�z�v���p��H�Q���\4�7��t`�g��<2�����z��6^�I�^��m�y9��8�P-à�2��ա0z��N���2�w��w㶏����z}΂m6
�)S���p�� #ql��,>�7Jbn�>d����m\ߋg�^� ��m'ޚ��5Y�2�l�S�Љr�DcJ�Ҧ�AY�6B=[��iW��z��N��q�n7�G{�
8}� V��Ѧ���Ѹ$�3�U�	u�T0�S����P1�=3����!���C(<�
����:㷞0�H�E�PZ6����I��i}��n�G�͒��_���@�v���^���;�~�Slk�n�BN��#��-�㜍�x+ħ�Y��I&��`�{r=
�����G��I�*�q�ɣe1����U��1+
XH��9)���'�奄eJ>��/�[񎼝�vb�"�M���Ub��펌�s.�"p'r���7�+(8b!�Aܑ�7��eV��q�21���.S%#���]�ے�ŧg�4�6���P����q��k`0�$��dB3�?;���)~��բ�����{��R�RX����eZ�蓫L(��w��9�q��JF[?6R���8Ջ�Tk��<bB����'P��-�@� �S�4`�Y��q3:��a3��iw���).�b�b��}�m9�Y�!�
�R"�����P0�6M�@�%�9���K��&�6 +����c��$1�찧2�W��~gvF�'H�U}z瞅:O"�p��U��b�'�Q>�|�a>��2`��Bh�\��Z����Q*�p��P�Z��']diΠ��H{�-Ic�������enyn�>bJ{�<�Nj?
�=�vu<$�m�'�f{w�!憋�eb%ķ=Սp��AFd�ZF�Y����8�����YU�k˖H9R�>�!=u��ɩ��ã?$���~��A�=�iQ�*�!h7>)Q�*U��ê5־�c�z<�<�0�7�#�4'7�r�&0R�܃����ҟ�K���|,#�� 1�$ü�G�Ic��N������7sn��f���԰X����{cW����@jow,Q7�R�с��&���n$�,~�������.�W �owJRj^�ޱY�*�䬿ai��-��Q��O|���:��sv�B��}�!t�H�����mt�4�d41Y]�5�:W�9�D�P�Jjq|� ����z ޥ/��q�kG��ih�	F�7�Mr�'���``uɢ�є��(O(�P��g��Rޱ����G�N�EtL�V5w� �B�0�+�2�����!�� aAJ߸П��?0������;4�4��s:_�C�@@�n��p��1N�����?���̴yc�M�fM���_��E|�#s��Ny	�+Ʒ}�.�C9��T{���Vϝ����h�l�q�|��6`�Ty�\i���Ѵ3H0����J��;T=9$f���l�`���F"k�@NY�C����}4Qt� ,uW�*�����a�-&ۥ7ע37h�
�IA�E��v�4a�Bu��:�F�3�NcT���~���-��������b��H��3�ѿ�\
j����b�����ir/:��p!��C�#��H#���KIA��Ai������Z�o��υ�)��@K-�q��x�k�-�IC�{�L�Z_�b�g;�k�м�
��q�,A�2�W�P�C7���>F@`��{��X^�Gõ�̣�+`"�CYx\�V��LK=���<"��������

I#�h��4�h�ҳ���P�L(z܅�΂fx%���l�,|G�*;ڜ'��k�j\�� �U�V�o4?���,��!Q59�yURo��S]v_>��j ���5�}u{���H�?�y�A�'�FGAep�7�Q:��k��]��	���C���:as}}%+#�,{�} �	7����RE��啗���47kz�3P4er�׏��'��̗�3^�o�W�w��$���,���m�������0 ��sI>�h���x�%)�gI��"��hR�ʡW����4�v�N����l�xb��d�6��a��z�qmq�=�d�}o䙏���n�Ӣ�љL��lH�U�͂�/Ģ`y�L\��X�?g�R�5�/Z���{i'p�����QD��%ðUȌ�&�J�ħ{q��%%�?�-TS�8g��y���f��\�(�@�j^�l�KL�u�T�Ɵ֔�5s5˖N�P���C�p�5j�T�~	#���s����iA��xxRɯd�bY.���T�er�d��S���Ax{#�赏�i9����G�&�м'FK�䅠S�oi�l�=��2���OE�H�N̉ܭ�r����v�`��������)��~��{�<�S��4��ty&'^�j�X���J���Jp�o0������o�����lX��>��A�5�b�"���zzŷF���E7������^����t�*������M�,�<2��6���%�V�*�7c�`�ے� 6���g�v7ĘZR�V���3�9@��p_>�����s/��HJ��w�\���g6s���������BݢS��tu"�}`���л�-F��Bnc�^O��>tk��Uc���c�d��%�bP��&F"-䅉^:j܋��]�H@yn����a��\�������-� ��M4?��\q}��::�j�v1Ij��k�ô<��)S%I���^�Ւ>t N�*ɹ�bFmo(�R3����ᕲ���l�#���CڟS�Q(&�%�z��~�khM���鐲US������:;�<������@�ߞ����Q0�nB9[^�^h���Y/�b7>�ҝ�ۋ��]�*)�G:�T�ڦc�s�S�Css��E;BpYs|��!'z{ �%�I���y�}ᇋl;����j~Q:��buZ#n)sT �����+�M�a_��"n����,�	T�ő�T�mT�̨+=���-.�Cy�����	MT��
NWx�
Р����dj�	7(����8������9����Vȩ`C��a_vD4o��C�Lu%<i��$�m�Xb���������FZ��lR76)�8+=���+b8Ƶ��Y<lq5+���0�T[I��Rꤗ�����r:���ס�{0t�[u���i'.Y�	�̄XBW��iV�Z�m�-�f������Gm�	E�>�#:;"8e�a��c�l�yk�v���	� �w��o�Of{ۮ��ws�@n��ä	�pM��9�W�e�L��9��<o��ɫ�������&wϧ�D�cvV"O��,�IA���n�D��Ӭ߿W�ǚz��hp�o�ڎ� i($/�H��p�����5T������f�{%:6�x&hiJ�R��&�2�w�Lv����̻�
���.����˖0�=���L c��u�ɋ_	�>nz���m��B��v�jQC�sC�v9���/CZc5�,��J��Y�>V�W4�y�)m����l�q1�^�u#EX[�%<t�'���&�}n��b2�/.��̄e��H��$� �;岎t׈y	,ԉE0ׄt9�F�����=>&�}#�\�|uQ�����L\q��N�~�YSY�n�D�1ói�[7?���D�6(�^��R	�6����0|��Kt��gwy��|�w�3�fJ�?�\hHe��ဆUR����u�xqbq[2o�%c�W��B�-��Y�s��
��8�r6��=�	��0�}��Q�(��y��ϖe�ڲS=$�O�Ųy�6r�2�����M�Z�(�͉<�TJX+}�k��pZ��,042��֏q�?�F������",�õ�w ���	�I��*c�r�N��N�j�jX3쌪���2ǌy�vZ���6�mҥ!��+\�z����߇��V��G��4 ��� =������J���T�/�OV:i��f��]M��
��ϐ���)�p�}dJ��8}�%�
�n_���M��u�5���3�������3���D�fؔ�r�t�E�xٯ�^�Y��\CT;N�MG��g�`|�0��^������l� x_E֍��/�ncOD�� d��1M�'����*���2t/]��G���Q�[���N�^5#J�G�$��3���v#a/�U��;�R����(4�%Yj�	��P�
R���.����D�F7%oL�4v�Q"ʦZS��l�mFg��G��.��.4:�S�u(� �~7��;��-�T��+d�\�!�9��c��ܟ��-�-\����]�G�G-���( Y����@&�i�(q)׽	��\��m�e��E�c��э0��A�O�g���4O/�7|][q���3u��sf��C��^养@�48�˟���]�`�m�I�0����+ɉ�l{=աd'�?~a��TFF�1�(vaLiN���T"|��� �i�dB>�8D�l�/UV� ��0@�#o�*�{�ˣ�Z�cl�r��r�"�cƁ��RM�bS3bV۪=b�ke�s���D��e�?��qY��^�OQs&5_�α��p<yC6!�9MHglG���^���A���~k��"�loKXq�
�e��fI���_��R/^�T��h�r�5��ϳ����!�+-L�Ke��m�ӓ�n�3D�ų�.�i�\�O���L��YmݰE�fR�ɔ>��̓�ț���o�h�=��������l`�t���~p&:]g��q2})vu�0�Q��?cr�x�Z�PIs�����1��1�_�Pn��S����R��f�����99���ҋԦ�;v�5��I�K|�8^5��������u�f!udD�rD�Hi8�-�.H3e'�]�,f/v�T��W����#�/Q�2G�;�7#���P�����у����q�C����m~� DL���yp`�%OC~�vo�`1'H��F������IG��R��t��ɠ6P��x[߰q��oHטC�I�ڄ4� ���Q�.b�_�,p ;�q��.�z��g:=��f�5a=���P��%5��N���r!�t���U�w@x3ƼՓ��.��lI���?A�a��;�	(L���ej�*e��{Y�P�ۙh�t�
��ѐ�B�Ϭ �i4����ji��9��Z��S��/$� <5��^��br�/�^���6�ή�`Vч8h���N	 @��>�sK����=O���5	�+K(��P�UJ˩�pE���>8���]vL�sGֽ�E{�Y�D��05`v�
�W���O�a�kpw?������K�9{͢�?� ��2&+5����鳪2�Z���Ҿ0��l$[�Oy��{`�ZO�d��!wGl2�x��x��yI�o}R�|8�[P�$�.�ټ�]0��І����ցI�eP7|M.� t �~>y'���{��`[x��i%��t�J�X#؏Y�� ��_��-��P>���p��$�@���J1>ƶ+����L�M" ~Mr�!.�9��j��#��~~Gi8�w/��/֥���B�x����I�Ó�+��G�Mޜ����;�ej�˼������V����\|E�)V��rC���Շ%�-������ȖuA݈_���ғjL�����X�/8we���2=ے�4/0=� �'�d'B��fG�彯M�k��Zc��#��qg��`Y7�;�y9?L�W�r��FN5(���b��y�e�]��p���S�lE��S*r��>�C����_�����)�	ċ�/P��S�7x��\if��s�ڌ�l�S-MB?5��)C�F�I�a�<Ўu<�z�W��Ɇ�t^z|����2�p�������K��W�-m)d��K�,b����En(U�>�56�Z]��0��?�&�!��3_� I����KK�'-NQ��ܕ��b��j�m���#Mf(�!�s�3ߟ�j�=���,9�m5b��fc����i��!' �}Q�����K�y���-@�=ɩ	3���GqM�������+���S`��m]���kl��ُ�F�� eD?x�5���7�sp2�Qb7T3U�H��~!)�w)*"҂�%���@��P�!�U�)X��
��:�Z��R16F��32�-�S�I8�/����\�UP���d��X^76�����QĠ�bEMf��V�k�>�
�R��x+X�@� �h����[�����$,�.�N_�lC�e��~|���J�^�������j�q*Q�'�ubP��[/����T�$���ʁ���Q��X�i`V\h�_V�<40Lm�)�#D�T{�NK�K���r�S/�dn/I�ʉZ��5��a>�ll�Y���m��Lc[z4��qf�7�i�=�kS�r !�'��k���>Y{
!-AR|"��³w�ۘ��9G~A�sKg�QD0%3��$���۔�wz�j�m�!�ɑ��?B������:�jAG2��H�q���,x�����y#�d
���p�tJ=�&���G����6�wx��wr�rid�G8��	�&*]�?�q�9�	h�wK��^�3uI��\Q���o�g9lύ��N�v'�E���`ӯa�	?5 ���^c��.K��)8ǺU'+U�����ѽ��b���V�b�B�����6"��.��:�ߕL`������v\������[f�KuQ�a}14���	Us�(��SN%�Sa*:�"p����uMvAC_DD3l
��B�&.�߳�S:	:��b~��K���,`ů���}Dӯ�@l��v?DYBǘ�� )�&~{��&Y��b%�����W�N�2Ύ�4�׉�A��9+�S���lu;�;�'>��cs������U�L���0�2�D-t�M�XX_��j�x�\R��
�{?%ti��
�_�E u�OɂF���~�ׁ�x˖i��Q�0�D#4ꍻ;�J8	oy�T��j:M2����߈U��ߧnc5a��g� (����c��?q׽�0���.�y��d�E�E�(j}���S$"�T��K�I��H��zS���h��u�N$�����9\Im�e�FF]3��h��ԉ(~��w^��ϛ���i��*0�����}[�Y����D{�Aɽ�ah�M����_]>�4�,��Ux|@�Z:��e(��V����R�VIzkpzgC�r]o�%���Pɉi����.ܟIb:`�� B��F��-nl�����r��W�ހd����D�EƷ�'w�����Z��5�ԓ�x�[�?�K�Jە�$�i�/28C�d2;ɿ�T�5���9C��a*u�F=����ŏ�����DX����:��C�5��&D�m��%�r�g�F(L�MEQ&MԿb��Qr�g�UO.�Ŋ]��չ�?�����'v��� ���81znJ�5艇�{ޓP�c�'hA(�<��JĎ��vǌ�1���&P���� $���$��Ob�K_T6+�;����y|�V��o�.�٧)�҇R=����i*� ��4�ر�?0s����=��%�P�����쾠_��~��w8��aǕuX�q��G�қ�=q�UfN��� 3|�4g?r��f'��ѯ� ,YR�������,q�Ȩ����
!0K�|@8��%�Mb �(�b>#����ID8/�B�%?-��x/����]��R�U.}�oF�:"耶o��C\e�YN9a��N�9���y�Yŭ�}LNo�ŇFG�]�3/C��|l����X�B���K�b,UuQR̒� <�p٘5I��4֙�Ww��'�wݠ;�o�8�1��)������d+����*C[���6R���'T<{I���xKX�Oy� i�HO���M~Ao���yBcy�0��"�.�+�l����:�4ԟ��+o����A��#��w��A�,��]��#��C�ß�hE��^6	M�]b��v<�r~u��m��k�C�ٱ���xs���!�s�.&��D�n�r�G���`;*�_o���;q�Hew��E	�D�o8��� �� �����@��M�K��"[�M�܄�F!K��M>�?�F$#�����@�M�Idx ��J��ԴM&n�qx�?�"�rv%�C������LU�4vcin���Oi�'Q*�J�zs\pF��C���m�D�����>��Z~�!\5��f��P�T���W������[ �2��j��X�\�	r�{Qg�w/o�� �:���;�>�D��3��*,q;��EA�1J�c�,̚�97a����
�:>+� �y�Qln���h-R��5��Gc�D*�+i����6ѢNdr�0�H��8���X�]���Y��L�H��=���Vc?��  ��:���&���Oa�/m��%x�E�]!�QU`"VW���#r�%�\=r��?�p�u!T�eҚ��zd����,��	�}�0���tc�"5�`����#����?��3a��#r6�T`�l?�P��$�S(a��]u�:���?���N�CX��l�����P��`����-/��Eh�p
Z���^W��P�1,�@r���q�绘����w��Sp��f��<��D�	�/,��t���-�I���Q,�5��q�n0 �@o.X���:��J��}�b�j~
��H�U@00TxwH��"+'����Ŀ�F�;iJ~����\��,iOS�ϻ�?n���-�Hz ����կ��H�c�i$�;���6� �t.73B��X2q�vbI��Zz蛚���B6C�����r�4���e�k�:m��D��u^>�Y>Gx���C1Y-*����jQ�*��
qv���q/#o�<��GFRI�����Qҭ��?����x2��i��y�oh��f�wSI�����Ӕ�y7�ל�}��4�"�Ŷ�\4+��$�[=:��Ø�^>zQ�E�z�)����V/���Y�;|�e60��횜�?�OU%�h4�
/Ŭ��GJbKXak~G�2>Ad��<�Q��}/�M�ӍbSH뫵�PҤQ�w7��;�!��#i�%rp$C�'�ӝoӄ}���\w%�(EuҌ��'I��Oz���>��lB0<sQ�����xc2��>f�.�e!�BQj+5��s0X*����U��U�	�U����B۫8��SFI:�������;����H��{��|�WJ��ۦ7�J���]J�՚���7j����e͗ ύ�l��8RΈ�q�f�`5U�4>�p���Y���=��]�с-^�ܦkUlrz�U�Zc�A꿒����^�W��̧�Q��cJ�]K��{��_���H��l��1T��z]���v� P�D�L��Jf�osZ"<�EA+W�'�c�ٕd����k%u�~������Q��8'y�OU�ګ_���-�+��!�+��j2��`�I�+��^��	J����������6���犚�f;D�~v�����S�-��C��b^!��B#c1!	��e����	��X-��ƅ���^�˪��ϗ��Ds6{k��Rt\5�LU{��U�ב�3�H�(���0b-�!�i�{�!L�+y�ɳ�����.��"H3e�8i������.�֒�WR���w>O�l_� ��p�X�%�;�dW��b����?���f_�����]D��Mݑ	��I?�	��:�����ϋ;���(abk��B��Z���57�kڸ��떷���A�#�b[�W�a�$p~�{����QE�.|.�ֆ ����y%œ�-/��+��x��l&�^���6���}+�d�Fs[��.�����0�\���$KsR�����!i:�˴F�����֯��?:T2��Wx��x��y[��lh���řҘ~6�7E�{�`:�?.-h�rg���g�7H(�q�Y"v dU;[
,$�_�3�.���	㙂7�P�s��O� �/�\�5���)`��99^K��1�R����[R֬jtɕ+��WLM��ڥ������Mb^~f�7C@
�����e7�&�6���F��.pf�%Z�_���LW��t����=�"+�{�<�	���Z����B̻�D���	N[����o[.'���r��(��"�ˡ�J��!����3�t�,�* �#��w�4Iu�"�&L��˻���}ǁb٩$Sk\5*˚�\��h������X8� �rx����Gd�pS�H+@�[����_M�~:�ބ��l��w��e��@�&Ҵ	q�����#űk�K���szLﳥNi�������>�Ҏ
I�fS@��Aͥx�PLx�����W�۔�+��:���c��!9H��%���y��ΎhQ�{��Uq/w�����/��W$�����o+0������c��UG,���eDg�Κ�A/�-΃��ՅeS�5 R�=�\����	��{���[!"�c�S�R��ѱ_���U�p�$�6�\
p��w#&T+t#�JP��L�0�F=7��@G�#��O�q�흊H8�r��֓|z<"�����q$�*b}�ekw���b8}Vt�V"�?�W��F�@w^�J�86�Ȭ{wվ~���sj��7��0��Y�&-r��in�%z������8%C�P*T�?��*��Q�e�-nP���>��\�'n.ʬ�rQ�Ϯ�qZlx%՚��-nĎB&����o��y���F%��B��O�v�!J��Ғ4�*]�;�Y�3"���&,�b,uJ
�CWŸ�����P� �&�>�h� e����qJ&��!��ro�4�~ӻD2a�iФړ����/ya����d��K\��h(J�Io���,@��j�����)�*�Z�CM|G���0��� �D ��Huo8�l����ʦ��^�������F{���l+����xH�+ϩ��c������[�<SEk�6s�?yl.w�I�&�ƑA"�2�}jq��_�}����r������I|�Tڋ�*�Y�*ͥ����S�Fm��R8!p�HOt&d��\1 Ï�L�gp��l�X����C{I�BC����iz���᳍h�{	%������!R�=��gT)R pF�noα�O0Ɂ�u@~F��>OD7Gwz�4�������u#�)�(���+�Q��r����v�z�_����?x[��O>�B6�H
�SC�(����JL0B+!�Ͷ� "���n���{ϗg�c�:t�@�-�4�n���;th��y����K�p`��I�T�c>"�������y�y������&i�y�%��Af���v����Y���a�d���N�����Wz^e%)�<�aaǙU4=�*�+�CYMgN�,��9�Xf<���䙫���̷�Y2i���{��o�}��X���ᘻM�V�%������15�W&�B�	���5�Ǚx� ��é��iٍ������W =�|.v�������B������8�V��C�w[�ڂ��q��k�y�ܟ�'��)=�r�$"�XC�{P�(�!�nIl���+���TĤ�G9��4,{���B;�K���2͑���b5�_�lp��V�f��������=:�%@�5�[{~��H�M���:��
� 
��c(0��D������Z������B�Qpz:��.ϳ���oB��\��Y�b�[	���.[9��p�;�,O�\�|P�ڲ�3o%�����7H^d��3�k�r��0Q������މ�o�7_�$��A�:/cj���Î�;�Rt�L����GF��s��>�\BCĄ#�h�m~��
^�[�c��f������q�f>F���Z>�d�
�Ez��K�ML��zZo��p��|u?�HV<��C�+������ma9��9��G~��t����p>��)�4q�Sr�z���� �%��?Gh5�86�@�%p�ֶZs��������~�$;�AL�C�v��ȱ�؎j����~o����5�?��Vd���� zY~�AF�$"ײ��0D�V��Ղ�c����������eX�ś��Uz$��<=9]�- �(e��."'�ž3pNUrQ�3*4��E��+�hp+!K[��,2"RL��'\\�
0�K�D�3J@j���\d����jn�*���@��Ϲ7�ӊh�`0V���{*�\&�#����u����kLW���uR����G�����yo-��<���p��zm	ِ� }� ^����b��L`+��T���Xػ�5mM�`:a:~����%�v=�g_�n����^x�<�*��h�:����33�)֢u;��!6<�yy:G�W������h#$����Ma�v�gv�wmO�j=p��Ϥ���t��!LkV"Z�Yݎ�+]c��Njd��Zb�b�q�t���C��[@�(?�t�_�~J�3���S��P��K�7��ܜ_i�k�m�/�7���~qQV��"Hf@�����h�b�[A�A�I4)�P�va�6oL�<C��nE���&�)�b�K/�����0��@7_���+o������K����~�̵搵RH�󓯘����є��@�����8u�q�7@���@2 vE���Ҟ��墰"=u?ν%Y�!,.D �B5�$;> m���u1Y��'Hh�_,�H�K栤�9lay5�y~����{e���a\D�-�i� �i����_�-���:,���SK�׵�C cL�h�*~�3@��+��B9�@<��\��O� �Dd	�kal��؀�QU�����\�	|���^
Bg3�~>h����F{�_ �1�:#�y��)+����i(o��&����7X�R���K#��,UĄ���\d{^�Y*J�(��X��t{E�S��Ds�t�GXCL��>�U�^��ɯ3���&�������yE<%:슁E��x���� 17�N�W���1C�[�z�F��JE��(<6�&�!O&z���A���X<�	^�%�٣:5��~"Di̇�?!P�P�q��ЍK�Pz�`�ʴ���U�rɓ��<ѡ�D�R�1�| ?rx<5K��N Y��-�T#��]�g��Э��b��x��e��1L�L�ޕ!t��S*'��<�����beڈai�Ӽ�Fݼ�a���_����J�/A�������*\���%hp�����e�+���T�0��~�U��Y7�l�Q�Tm�=�_�UX_�/>D�V�Y��nE]�U����F�c�z����Iנc$�ĭJ��/���ڇd���3U0 ]dCr�đ�*�<f�m���� <���=�0ښ5 �#W���%0qD���4窖}tԹ�3sv9��z�6�#7�^�ƒ���x�%L:���A�%V�!=G�'g~��ւ}���B�?���S���-/d?BU*D6��<W�|,1`"�,�3���f�H�g±���00Ѧ��f,�l�@�摎���{+6E��+���Ρ0^�Qt_e��f�VG����N8���Ʋ��X4P��G���PܳI�[����>�,��)�cN$ԁ��O�1d�����ǭ�QV�D8d�4��
&�*��B5g{���C"�Ou�`}'�Ќ�62N��,?�'��hH�l�weXt��g ��);��G�5����@�G�L�F�8����h���x��Yr�EԒ��æإD$�v�.Zy,���N�~����Z�TY�O�	��E�ko���ic�'�˞��fe3�3r^� �vn��ϡ���	Q?��Zx�x*��;�M鑰u��.�TAT�r<T��Y}� �3&.\�YXwo�a���X��z�R�K'�2�OfзX�h�dO��A5����� �f���(i�u�G�j�������A,��#�Xvk�x�1�=r^ȉ�0_W I�~O�>p���^����*x6�^�5�ʳ���������%|����[,���۵�!�{�V�Xؔ0��N:�[ǳ�f��څ)��n 6�ea6�Pf<a֓p�O}�W�7��}��TN��}��c�s���y��޼{c2���A|:�ܓ/(������qSӰA[�y��2��r�r�;��W)b4)3g���9�ޥ@G��6d�ī4��Ӵ�ys�heO!s�F����GY��{�uk�KMH��Ս����?��S�d��POetͫ%� ���4�Q$�"G�K�KU�v�%��v��S.7�_�B@�T�� �%M���b������j� ����<��VL�[���k{��hmҬ�g���,���]��-cN"Ȫi��1
�j_v36TO��~��&i%�_mψ԰!��,)U�v��z�����r-^��Ř�}��D�+0	*i�m�-ut����������rd�3s�D��b�FW�΋fb�g|��^��ZwkTk��W-/���޺��O�d�y���QM�S6�5�E�]�Dz��T��3 b��q� y�e�M��G��V|"�E��M����M&����OL < �i=^���;�ʆ�z0�r ��6���5������Y���uC�n�R���}�D��kՇ����2���Gd*g`�8��l�yR�+BE\2���a�(��]��>�:��(����P��	&{;tA�J[�Aq܆�ݗ�9LZJ�&RT����(�3q	��B�ُڇ�6HI�d��33��.��4�H�����=�m�z��zd���ӝu�?:Jx�jLP�|C�΍��e�%J�K��[x�ʍ�oݮ�^rb�O_�堰<��C�6��Rm��g&b�0"���ch�4/�Rc�P�V������H��?�De��{����+�-� ��g���P���@{��jv�̡!�`�R�Q7FT��B��Va�BK7����ӭ������u1k��42�Ȃ@�.��C&�u�5�Zi����8VoG��Fd���gO����ɻMx��C�pp�x	�ɬm3E,�����I(�a�=����/���N�~T&+�C��)�Cy�T��2�{{NV^��1���wa��)�3��\IT��j	�KM�8��&P�ӑ�/$*�/�=���m#�/D �C�7�iD�cF������V�"WڊD�ű_VMa	�(6佀��VGW����O�r��be�:TUJ��b�AMN��>�w�|U5��7Ί��l>�Q���{�goq�zE��'�[�Õ��3�}��k��;H�ة|��)�5���S����)��<�T�MLXJ�Eڐ���)�r� o�݌��✈a��:M��33�&9��Ҡ����P�%	=��3�4�������� �F�Z<�	$�WS���Zo�@q�wk@��+AgEh2O`y�9�^��5t��!��C{��4��	K�P9?���_��I\��o�M�"��x�5�A[��8�reM@ON�nav�P�^"�K�I��;8h7���k�f���DmX�yzH�fc+E��2Wq����єBVQ�����/� �>��S�*�(�#pO������=	`w4��<a�5��Slݣs��A��+V���������TH��T{��}�xg�ol���%GM�8x�d����C%>b6�6P*X���/C@Ri�r�$�b�-���,T|~,W�����j�%TR�R_O�O�)E�e
�!j����&2��#�����C��m�5�/9�&@`�l|�g�B�����D!�@|q�����6Ŗ�c�k}�ß��л��靮e ��*�wٽ>�"��c����7��ri����l7s��6���.��@����J�q���v��H���d�3O3;]hq���]	T���Q?cvk��7��[%�?Q��E�9A�T��V����D�i�/ o�%T�woVW	�y�.b'2Ia�R���,g���R����i����C5�N�t��L���U��5��v���-������rڏ�c��U@v�/���ܷ̪�e�w���>���M� ���*[0.`����vXc����g���>Zl,�MN%�t9\D�~�Ip7U�V�9�g��y#�Ѷ�f%K�|۲!m�k[O�����B%%=��Q�6�=���Ke����?��;c�׃j�_"�p��ͫ�z�f�ޟ���f��#���ٛ�$�9�r�-	oN,�f z}Q��陦,��Fބw@'����w[8�eE�����{�vq5��Mg#2�/"��/E #B�܌9�aqC�?���v�rq��������|ǥyu�*���f�˞�U*J��LÉi��+�'ߥ����v�R�m @H �+��.�"i�K���[���E��|�������"W��Y3��C��%�R	��L��$����|Hc��a)�:�Hd(3�tjO��s�����6G߹Qipb\��C�؊�
�-n�_@��=_@&ZYJv����IxC�Q�7Y͇z�|ݜU��	��9n��G-�6,���1.��N`wg�x;�u�̖��vN�Ӛ�V'g�o=���R:��g�d�G`�Hjs~�a0������@$e��*������آh��qN��ri�����4ۢ��j�����GA�׋�5��&��V�OF�]f�\^��#;���ں��!Q���ቂu���C�o����"��@͛���'N�\>V�;vE��5`F<ǡe�A�}q|��L\�0u4o��D���b��_ށ$�>�#>����G�+���$f�?�&��P4��f��˰pa�����H�?>M]8F� !l�.U���+���0	�98�)�d��~x���/ ����bk=��1�% &����vz(�&Y�1˥k<��D�#�(�jz��*�l��q���͋ԅn���R�W ���/�G�
�}Ђ�'"͜�Zm�y��>����"���k�b$��!m�U�
�>�N`��t�jL<R��6��9��n������'1�b�,�]X���;(�M�nrg[�q->�I�:�K��Xw��՚��B��Y�"�������1x ���� �=����n�
j�S���tV+fq�h��o�L�IOЊ� 1�\M�� +�@^��02AZ��ǉ'��z2u1�zk(��	q�G�!u��o�T�.�X4?om��ڭ���Dx��$����ٸw3���y:&�D�Ptɼ�`(8�j���-���ٱ�Φ"ꌚB}���v�z�.���D�?Y�o	��6��;�[*�5���	HOOj�M޵oE{�.�x��W5Ç�(ګ�Z=�=oė���� X�)��4 L1,�t	�2�ib�q����X�9"Z󻄏� �R�<�4���@��g\�'�{ڢqx<��fׄN9�Lg7=�jgd��B�b7�"V鉻�4���$c�=�{��ϲ��z��YԤW��"���gp�c�]�;�R�2�/���?��izXh�:���MJx0d���}��{@~��pq>MQ�l�Pg��na�M�����*H؟f��s����J�a����A�>� c��_H�9��st�F�T*��W��@O��G'�?܇�\�VJ~}���	�K%���0D������[q��`4b�iX�u_�ӗ�����_��R��
ؽq�Le�G��ZQ��� �qX���>�N5�(�+�S����:��20�Bb��$�6�^E�x����O[�
L(60�B���9��zQ����_��@�g��2N͔�'0ZЯ����i�J\��f��id}N�gYsİ��&�p�qn�I����U!�<l�J{KI�Ƭ���v���u�o3H�@eR.�X?��?�՚ҏcW�i(3�-�]�2�n�E�%c\��-��4�]����>��0bt=�����F\oa�{\8@��Ym�_��smk+���`n��j�yk��e_M�ҙ���1����21&*�6�\��`����8��U�����S,�/����/�Fr���"���j(;ZA6IӚṻ���hdb��O�R)^����Ж!�=��E���Mq����}��3k�ڷ�79��:�m�8<�M�[wK`�BQ6�| ����R]_���C���8���E#+����_�SJ�pQ<EM��{��v�юlQ�CQs6Rl����%G��-���к�H�n�.�0�1I��`���r�E�t��d�������S���d�zN	Fcl%n�J^���:a6��%!�����F<��6�*� e��}C%D��\�������dz��5Y �!T%jR}|S����Ά<��B������q�>sh��/բw�b��U�b0֛La�sT���% T���$��{G�q5��A����?��t� ά�݆�<)*�{Is���Jh��is<N�/�K��k����>�*�W��.q��.�c<��Ӝ}`F�X��1v�['��w���K#�o���-W��T{��]��l�L$�eTD����x���*��i,�_#�Z:��F?/A@�aR'U�ĵ�7.C�����Rt֥�L@3���z�-�l�9^4o�>����4�]��㷱v��ڳ�I���1��� O���Y�
`�kC�F�E�H�ic̀��/�3rPi��{�t�[Q��t��KO��E�8w��C�~~7�D?���ay�`-x�a(嬫Js��jKMy� ����>�0�D�.�P�(̰�����^�B�5�)�0znl�����QãLӦa�>�����7�f[�!L=G�\B>{��+�;��8	.��HX#<�l�z�a�/�..�]��h1��ppz�w�q�L�:����pT�Xy�kW&/'=��p��4�� �	��(�K�o�a��*���=e=s��Tٔ.4��;S^9לz����8�������^h��Y�9�_�w�!�۵�Bw��#>��U���tzf�I��Cw�G{*����~-�n�AU�����Lq;�Ցo�(Б��H!��]��ߒ.��r_)�)1$�D��d��@p&�XSҪ��[ဎiVZ`��H�+,Ji��!��k9r;��َ��Oa�\���~ZR`�qa-���Ϣ�p$�g�2I�f ��f!u���w����HA)������$r���_W��`y�5������D�X3�=��Z.��;������_��q�h��~ /H�f"�fv�T8�z]=s� T%��wɤ�O��$�J*
��[��� �iM*�2f#wXA�����8����Y�}<������Ň�/�` �K_���ϴ�e�ؚ�9�P"�5Ox���-$�1�W/{��^@t��.LPD��w�-���bdt�R$�P�ڈUD�K�@���K��yN%��7,���aL6E!�*mR8*Q 7��Q���ǅ�<��=]F�=|�4�b�I2�	S� �~�q�!��a�*�?��ޟ����V�/�V�7��q�����^=�A'B/���3q'>��l��x�>y��6t�ǈÝy`�p�"%�6[���3E�{:���Ed�AW8�E��b{_+�����4ٔ�o&(��P.�@�"��/�O��B�33��7�h`��v9�b�`����t�?��D���^��ہ��-�0��Ar�b�cm&v��J�Z�����S*�)n�w�7̐i��P���h�JH�S��rPX)dY����.�R6�u���xu`6#y@���\l�2jƺ(,oi�24�/u��;�HN�F�������������%W"�}�K)����;��gʂ-vw��Q/z+�[�"%ߖ��O�؂&Vf�n�l��z�K����1�������&�@vh�@v��cw)�Bo��K6`��ݡPs���b�J��k|񍔟.D�Э��ʨ�n�h�]����Μt<�Ho�}㉐c������]9j��w%��C_��Y*�	<���Ᾱ��-�/zZ����k�}��%�b�8���:26?���y6C�7>�Z]a]񚏫4YP��#2Z=�؉�P�$ɂ v��+�lAs���H^��~�|�/����i���7���n�U�������/�o�@�m����Z�᠕�3x�?5�ט�����)���g��ܲܺ�Rc!��0j�����^.��*�w0lQU�۾�]�px~ߴ��&h�L��l&�=��fn�㲓yǯ����e���6ߠ���
X����4�+�S��#AE���)��P�(�\-V����7e)mE�-%���:F���R<`�~����L���e�7J��YR�S�Y*иv{�� f}?m`|��v�z]1��N�,��*#�gP�Wy�ǡ Pr�:~�yߙHG#�dtT˒s��^��'��������U4������ɽ�יYr�H )�佋��`o��,:�΁5+:�c�(M$E?2�!���Ǹ�o�lq�r5��o����V�?�5�M*h����ciA0� �2�!@DÉ�Ï���嗔NR'�� ��mj�_���^ ɽˍ9�Z+�Ѕj���5�"��\׆:�I��<)�]��a�u�zhEM�;��ltJ�B�Z��l���-�˝�r��ٖ�P�$N��R1T�Ҋy&�/'`����[}�����龴�9İ��$;t&Q�H�Q�=lt���,w�h�R<�K�%M>b_�Ѹ�磿8��R���<�\u���P�_O�Q�d~ `�֪�ePn�c[~��(�q�C��OS�wDuU��"1� ?�\z��/�П·���+�b�#k�`�,2D7-�c{�ωΈ��cv��j-�E/�S���-�I�t�}�N62��Dzh�fB�;4L����xZ���
)ICϔ�9�¥	�RՂwM3�E��oȑ�@�L���>�G�Kv+Eb��b��7�m�3�wl��������jy�?������_O�*L�~��m�s�H���	.�[9���!	��~hh�D��B�b�N���\��ϲޢ٢�~WP�G�y�=/wTV�o����D�H1��F���$Xbˎ�^OhޕdqQ抇D�;.�c֤T��̍fj�e��u�mv�o�ʍ!{��V/uaìLJ���Re��'�6l�%=M�ϣ�����m8[C�(I�y��m�o��֭\@�K�4��%4���ǔ�<�B�I�=u�C�"��M�E�P�L�~�t�}�Zw���X�wwg��u��q<�ېY�e���|(.'I29k���
��b��������4�)��@e�i������W�o7��X�S mJ[�e������a�^���*/}�������
�0����9Zs.%@5���v�I��v���>8�v����]`D��K����%�"�<�!��qbdp�j��|Pd��c$��B�m��tA+9�Z�|�Or��c@a���/f�y�5�`���o/�������V�Arh��<��#I<��%� ��x�e����vR�ەc�#rOO<���>���t��q��#H`ň�*|B#]�G�JiS�U����B��e�bu�y�6�G��o�5~R��b�t�?lK��֪ɾ�e꿿`�F��MN�]U�?=�=?xX��P��3X�&��y���RQ�=^<�ю�I���+��O'��܍tHjD�� HQ��Z�H�−� �-������za3�ǖ�nF��E�y�j���(6��u˫�g_��=D̸��l��g�5�BS��1,��w=> �[�j��3_��HR�C�e%�[ z���EE��d�0<8Z��ۅ�.��X���ѓC��~C <�Xy��O���/N������9?��௉��Hz�.7�?���ZritD�/�����םt����0&�+���^:^�9��0$��ۨ��l�n4~De�o	u��ْ�q��A���R��%�j�G-ђ�wK^Z3_��٠|<�=�|zE�h
,�R=��A��d�F��Z������f��Ȉ�G��1��elC�$g侮^pR��'U9��1gjS�FMR�I=g�H]^���y,� vg�iO�E8)�ET9�Gыwc�`5�O,n��VB't>T�^Q� �^�l0�4�h��+��n�H�����4f3a=�%�(Щ_N6-�M �6
7��.؀�l�ʶL�Q�	�Tr��O�{yra�TH��O�z4���A�s�'�	,�����BB'�{WG�薮"&�]3^��yz%&��(��˱9�)�߮v��w�z_�����9&f�Cp5��)�YTƣ�Pd� �'��Z ���P�m{��Xըs�����LGFB4��a��I�����c0�է7��Нv���A9M2ۏa���@�n����umb->^1�5��{����ܼ#e����Z2�Bfz���ǝ�D8 :�T@��,Ѣg<����f%�"�t�=�%�.����%�4b��ܲ�!H45T�K��ؚ�:�9&?��B:���l+D�?�κf�>>�<(�`mS[B�O}g2�tA��p�a��������v�M_
'�'��Wdb�۽��y5?}���vg9;e-����ʦvG-��xs����ԝ�}��g�w��e�9X82<V���j�_������e˳þ�+�چw��h�	_��W� ��9}Y��ÿ�o@�N=*$��0�1gC:�T]�de��ԅ�\�b#v�52�'N��7��� �49b ���W$�e�̬Z��*�x�j/֞4/�%�;}��~1�U�\�Q�5x%�)�=[J��X��i�-2z3h{n��8�5�Ҧ�fy�T��vzO{�܊ťJ<t�bU��&�������$,��L�k���"2�����R�#.Efbn�5#dƖhE��Tl�;29hW�0&��k�{ �L����Ò2G��V�C+��
�4�@�A�gF}E�x�H��W-9������`�|1㞂�o�Y�T�{f�O�z$����;$���)��$��7o��rx��
 Qiy��� �n�]l��D��%yq}���n7�p-@�C����e�ں��j�Tr�_}�8G�������k���8|����3�SAcY��%�@�̽3M%V��c`�9̯���\$c�|�h�#ao�ODE�Q���ø��xv�@��X�#;��{�XD�$�)��kD���_�oi��'�*_�� �	=��SꧻlT��Gm7wcAJ��j��?�S�O{)�NoV�
=n�-a[����D2}4���x5LZ�w}�1��������h����^�iq���8hU[�DH'�3�_���l�p�����b|�zPA�f�f�G���G/�+�VW��(�?�2��避�������]-��a����݃x��kJ�Z�����?����6P�F��bV� �p����|�/d���H������'���q9Z������B�HY4�����!&�D���Jٱ�rX1^�#��m;�������m'�NL�M���������ti~�PY<�	��󼥌�(m��S[�o��:,7wb٢���zJ,�D������xZs01�1P)�=#������L]�.�����`/l6�-U�)oi����]^\٪fi��jSv��^���$�8���uZ�긃��^,�\�c/s�б��i�����.UkB�eO�~,H������ԾՁ�y�lh�iކ=΃��e��y&.����^�n;:/7��/8|�_uY�S��t��&�꼏��p?C�IE���7J���{u���;#1?�%������{�Ev�����EzO�9����b�7�ҭ��N׵g@f�X9^��¸���J�5��}���pi��w|�8��K���2���v� yjgL�kI�N�/<V�����np� nHf�=�?�]rO����ҟ�7�^f�Y��F���h����R6r�5~�V~$:Fg%� @H���ى�kh]�dib��y:�Y��L馞$������	�F�ƭ�F�C�ዃy��*͂�;~	o<U������dv^�K��xA��>c|+Ä�<��.l^j��/�#a�_$�H�eZP`Qqj6��	U���p�L���a9V�v��ۈN��F[�!���#P�mg�t�~���*\�q��4o�3�b����km�␰.y�S��f2���_�4p�b/�b?�e1m�s��.¼��?��r�)v ˋK����v<#����.1��#$�N��OTƛS^Oʃ��m�G�7������㌖�j3h�ac��P���7�+RO���~(Gy#X�v%q�_�����c^�w�gῷ�t�ߢ�?؄�n�S"�R4T�F�%I���u�����i���%W�. }���Xk���<
��������-�D���g�8j��2Γ
T#����#�T#�B�[���f�<��ZQ�ά�����*S�'����Y��K�3���!���`��4��%԰�\����Çm����1/Rس�1���^��6�)
�@���0H>X:?�b;h���7�j���u�W���+
_�G��M�)_�ŶCW"�c���^��(��0SL�ԯ�R1�Yl؋��V��y�6�U�)&��>O�М:4�-��2M��ck3��y^�Ҏ��[��5-.Z<�l�Q+��8��۹o�C��5��+%� ,��&��s�Kf�^B�&���qʪ�ǝDu�&fw�
���N9�'�ꣂ;9���Y�74��\�e}�}g��O+Q]�?��˅�1���1�h�u[G>�ܐ��]WΜ�ȹ��0�Z	�k�vT�Vyy�'܃�}d|M�荪.E���f�X�u�O���Z�[mHU�@Lu��mz �2��45��XӊFA�l�l�����F��+RM�0>rGA�{ ��N.T��^DWTAc	�xր�pC]4װ�rqAz�	ll>�&C2��ȟ��`!�Ngˌ���l��𯗻.+Wn�:���z���uu���{��tt@�K<L��6l��]���e֞��e]l�+vi�/�A�o�����eĨ���7��K�0����/�� T�D\�����Y����B؜���ZǄ�S��mS�:��%L.��_�)�' *�Rz�!��3�_�7�v��\}&P'G*:�81�ɝ���8<_ٱ~��~���P3H�� ��;W��Wi"!�&���Uh#e�ٮ��O8<h�t���V[v�_Y�}w��z!�{Z����a�b�%��� G�x�C��8��Gw��Ce-�K*���W���X={�٪�J�ۥZwJ���0B �x����q��!�l�T���U�}%�w�;�Eab3�f�聯�~p�m�����m4��?O��;�@�B�oc�ŝ���Yr��]z�iA�v�������D'��X99��v��q`p�'�!j��ui�D+Hv"�o}���G��8�a�|H������ʲY1M�	>L65���������12����O��/)�вAIn�y.^����bG ��p�
rv�Y�6�9K�����7 {9T}���#IP}WW3E��X��v)��^�jk�LF���2�����d>?�w|�����ʆ#x`��ʻ3#qK����NV�B�=�Uߐ����l�����:����B�Q�N��Qƭ�݁l�_��RD�BHÓT�]��ך� �qV�nJ�i+���b�+K�w�x���&�'kg��$m�N��^�hl�;�{��� ��'�#�0��p�Z�<w�1Q��Ϫ�4����0[��>�_)�h۹ߠx����;n�Qq2#V��Ya�Ղ��-�;*�d��	�kx�B:J,QP�%�A�\��V6$�7�!��5����O>ş�/�T��(a���RiWq��'g�7��<���i?�>p�"���[��V%��P��)낣=����5%ڢ��]RR��1�]9��4������`��Gq3�:��E@�l����ҹWi��`��xnL������g��&9�]�L�=��Jj�W���xho1��s̱�N����1�)ih�T�$k�j�u��W4�3m�(���b�"��z�}-j���+!�o������D�n�)�]�+�aͶ^J��Z���E��$ʌ:�l*1�2��/�L�<���"{�N�Yǎ����\ˏa�^8M��8�T�@b���C����m!R܃�1�:�პ�Bd�8��s��)f*\�V?1������>V���M$X�KB�;rI�Yr�~ |G�N�Q�*�ĠZJS$"�%�Φ��L%�I���ޏ c5f��'�'�r���7�1D�d��((p�����*"��]�z�e���}ԏig4���}Ll3�B��+���A$���5�H�9�����]𺳾� -�]/�r��OR�]��9@#���*�tR�i���QIw�l�_����B��*�xXxw��%Y�X�{۟O��M �V�/A6�do��[��q�U�����=u�wK���S�� �A��/�c�]����d� TR���C��K�q��a��m1����GiM5TC�bZv��aV]a* \e�&mP��_����pM��	�\�u��� ��0;��bȭ���zǫM��t@C�j�?�mk��*'޳��Ɉ9�� ��5;��T��V�>��$O����g�aOS����
�[�Ɂ��b��I!	!9��琤	/��.ڵ|(S|��+=�����V�?�(�Ω	��O����3��;	��hEǪxo"g���ܒ�r�y����o[,�B:?�wŒ��pY7;:��b�곯�r0SF�@�WC4�CHi[*N�������=�!�I�h��*y���V���\����Lg,�J�#��O�fb��@��A�F�i���E�5���%%�k��/*�+��_}��r1�iq#�6!�E���Y ���e%��Ϛ��^��F�e�	&�,��ߪ��E���¿�X�:߲m�`^�d�m���H��d�-}o�D�Eo/�_�#��	�Ow $��H���84m�D}EQ�4x�6��Batc��%i��4�ߍ)�+�@�Py``0y�~�84ܛ9�bO�o%��Om=f��$�^%04}�ζ�6�� �,�h��!N��Ӵ�`z����O�[>�U\�yA�t�r�����H�Cr��qj���M�L0d9umx����x����:Ī��}��Yޗ�/k6�S�����=�>Lu����bs����5Yj/0C	m���z9v�.��cW�-�y�n2rmC��L�wl�@[�G�����ψ7��-7z�E<$����3�K�0e谲�'\զ��5��V��Na��0���Pi�V��K�r:S$1��'�@<��f���T��q?U\�խA��)^�=��6�F-�C�s�@Wf4Jh�g�x:I	�TL�T���륾�ب�\?����sꚚ�����Y`^mq$!=��9nA���׼�]�O�z��`�����tpت߷?v�i���� �^띚,��7n���JE?I��$� �*HV ��|�+4z"&��R��)�|�2����>��қ�o1Θ���oO�}��_��{��e� ��ԍ�C�%+4��D����V����ڂ)��sk|�I�!�G���ӽ�5�ݫ�f���O�����S]聮6�����܈���-�<q�;Kq C���Nn�R~`�3���	��:�aQ(˫�&0�t�=�bH-��PBNfS�-�s\û�B��K�r��@:hZYL�+[����t��K�$V0g�d��5����h~�2��~�
��RɠP5аu������ ��}O�1�3���ꓕO�K:�a��a���:�̙*��<�EG�}�H퀪!'M��[��������jmD��'�pF�P�5����n�kP��ݽ4����e�y��@��+�mw�j�l��ȳ��VUz@�VQM��}���#�%�<��Q�pM<�n�[X�G�����K6�f�2�+n}3�W/@q6C�W�]d �7��O��d�i���ʿ��x�/�Cj`�E6!�e�QNK���e�w�K8}l�J/H��O ��hꆆ���&�.���
w�fڵ�Wr/� �@H��xK	�>8W���~\y[�e�v(�*U����ҟ��N��0Usk4#��w�a�-R�C*0�u��9V�Vh�i�׼�K��V���Xq=��| ;t;A�?�3�u=���焮ze ���H���O̗�Y�nr0b+ ��GGq�*���v�X�{�ں뺚K����-��'��ufC��t�a�ۄӯ@%��@��]}w��<�L��͈��I�*L����݀��!(�|��A%��W�����V�?��q�K�Y/�;�^�NA@ޟA-�ȑ�},�p���d����[JY~�9�0� 0�{��h�P0��ND -E!k[:9�3e�8�ճ��|���FP\��oE�0���_HS�N���b�чN��p҅�4�akj�@���1q�:J/c��2��V`C�B�(õM��Ux}*�C�A�ML^ٸ� qZ;�y��w$�C��;�(		PC��I��r��&���I<~4�9W�vbʤ򂁋���`ex�^qCz?�?T��*���^���.?�����\�'e��U0Fz	�ȎB���~��2gsOQ�h�U�e��i�_?)��`ns��]d�Py��+�)�zf1���\s��$�3;�F����T�7�Re/E�2�:!�SW��|e+|r����~l0j)N�l�J~�~�%� �36p��X��ɫ���0J���ư$%��|u�l܅����b)9�@�I�:�����G/�G1 k��L�+�+����W^���)JRR�h�?���0R���t���	��	5f[��L�$<�$��r-�������rE� ��{'����MI�t�����l8� � &�Ͷ��~0��F]oH���S��G���g��{�E��M�w�7��O��28��>�n��i��g�Q���z,�@���ը���f<�gr|�a�=9�qN��n@�/��lƐa-��I�ڒTҡ��6rL�[cO�F�R���U�&su�e�h͹7�V�?�i�a�d�����H5)��@c�ܘ�0�ĶW��km���0�� �!��m��@��Y�8� 䳢&dO�b)��?ˠ��y.��a,�H�[����_I'�R\p)�K�o2kI� ��i" r
���p1MN5nߢ����3��`�v^�v��.R��4�`�����^p�"����H�Ac���M������p=���?d,�=I���򑊖R����[�"�y����g��Vkx�\��K�O�����%���N'jJ��r=��#�-cSV���_�-�6��q֛���1�NJB�o�Ƕ��9�V��`B�t��P�8�34
��q���)`G��$<��V��r{�J\�1�bh��V��,/N�x��F����~�+���t�>d"V q�q*N�(R*�	�Q���V��)���9�k8y��i{[i��b��Btik�Ր�,v���&�gBQ�L"�b�3O͎�*!��g"A&��)���?�kS��Dn~y[;�Y���}�gؔ���.��
Љ����������:����~����Þk+�m,�6z��sV�XG�S/W����k��o=��O�
f��$����a�_r�x��In�\�-��W%ҹ�K���lo�9K���_�uI/��]��l�C����W7�'#U��9%��xL�~�ݿ�Pu\�!W�B������z�D,�8"n�V�h{o��qo��#?���y��,��_�z��Cqqܡr��,��x�@��!��]@x�R�_�����q��x��7Sʎy7y�:���a������3i�����W���E?F��`�"KV+a'��Y."y%;"1�o�)qʦ��2�SL�d���Q�q|���������%x�]��êT͗�a�����7u,�}5����c��|b�����f�v�L�A58��r�F�Xa{�w�=ަ"�͜gDC��67�2r�RIn�9�1g�E�Q��(����)l͛cM�H%�\g�VnU/$(�:��Ϡa+<���x|��ƿ(v�k�XcE&��EnU�5��^�=����>D�Q�b_扫�pF֪N�&��� v*��@L��������k{N�F᭪��Ē��RT��4˽u��o��#'�Y������f͠�$�9���M�D�YJ��d����؍lV�G�]�9P�c4&(�5ue8��Ћ�f3ϔ�v���=A�Y��B~߫�����ҜG��(=����!y��z��<�p�:پv4��}6p1-��Do*�o�t�g_4�;�נ��D�g �e��+��?B�6V|�&�GTe��bL�o�}c�.�����T�!x��镙C��(( �~e�����bU$#��@�Y������(e���PF�Ew"v�'�N�z�B�Y� �fJe~���.��"�08m�ҎF}��e��Nб�rJջ
�0���9%,�O�-k*l��Y���c��̓��CM� q��:	zZ�@��?����Ж��w��P���r�5[�nc��/n���;��d��\�(hzn'��O��ݩÐ �t>�9a|�6��JgŊ���Xf�\����6��pN��� ���	��ui_�z�2c�۞}�>��c���^���7�n�L�`�wL��e]of+�<��m�^�C����6�������]g��T��T	��������[�W��e���+��>ܝ�$���:2�Al��ZFm��욎�gA8!0��x��5�Ȯ��}�T�i,?��0�Z
5+��b[����(�M�1Rz�Y��o\��LP��	foϤ���`ɻpt��t��R��[M-��}P�תD�Z�zM(���ze�:S���I:�m�����,��*!���A��w	-��?}�8�1�5f���ӝɟ����ʻ!t�d5U�Fi�ZjH��lR	�Z�*��d�)�̛�����A�u���<,P>/@岜�^e��Q�WZ������ Qbmvu-A_�->�^B�x�����G�^/|A���k]l-R�@�q��Ék�JLG"�+�D~Z-fK]�ԏ� 7(�Q��؉L�,� ��/k/~���K�a%�k;j��3;�1<2�
]��'�z���햝�G�-��@��!���F���w��Ǜ�k�k��] I$��	׊�A�n����W)����0LZ뻥��9� xU>�3�f3!��0ߓ2�/�8�1�����Y�n�/��/s�*���'z�M��S���ܚ~H��^a�~��,G��<�*ٶ��|�E��fW�SX־L�WvG�:�ˡ�z,����a�\'>%<�.�x;������_���\1T�4y�)���0´Z���RX��4yqD�*$�>,�qr�qCL�������đp?gB�I����F�zr$.�g�X�~�	�@�	 L>���}g��hl��N���ft��!<�����룭rCjd@I/�sF)?%O�FhRO�35�DZ��gt�F/�.z6��Rv�Ӝh�)!�p�J�yk�
��h݊�R��E�Jm��q�6��_�* J�f����*1ѡ�O���f!J�	Dv!w��z*���ܐ�(�F֏��Vӷ|��� �RS��r�{�(x&����u�Dw�=;�BЯ��H�&��,r+>�~׌�����'Ѹ�*�-�"����D�	�D�����D�����
���B��BE�����w���=�7gU��]F\�c��7d�.k��7�N�!�9\���Sg!$�%G.�Ϥ|�:�j=

���t�BЫ�Ƈ���^y[N��s�Y��Ny}$�}���M�i
�fy��C &(��$�x|cu�Eh�����Th�a����y�ˑUi�v�ߧ�� p��eUE:����l��8�5��~T6V<�]�f%�7*�l$�;�����z�E��p%K��Jn����q�x�Y&@�i�j�D6={���{�b�����V �VU�� 1䉯�!��G��x�*�͠gǛ���Aң��(hE��y�v�W��L�m� ���%�Z,p�jcyYޓ>���/(�?�]�^KЛ����5^Sӹ��ە�������F�~?s���ڵ��zw��V�
�����G�u��u��]=�5��rMd-"�%��U)�	�����O�	4"#iN,Z�������������)��:L�AR�����&,����Cg����!^p]Ko�3��m�E���J�ExguY�ԭ�9}��P'�@�Is��
>�E�b��E<�S��"H.���L�3�Y���׉a"���&��e��R��[�����{� a��Y�ĳ��0�ƙ��+Q��$�N۬���g�)��b.�'V
�^`����Qu�Vy{���5�֨�P�;�+�:��cc��� �G\CB�&B�:7�*k��T�_�/C-f�1M�f�=p��JzF^+\2���)�^I��F?�EzL��ɉq1�a�H��?v�F�8ZE�\)���},w1�k�a�nP�]� ��Cx,f;�P0=|�n���ݿ� ���m��:�9�%�\�� E��Z�T��S]St�X��pݷe哣�2Z)v�ЈME^d�7�?܍&+��[��҅5�KG�d�\xV3�1+D��KU+���3� �����J��.v�9Pu�6�1�G�͋c�y5ߦ-"?��w��I]$���C���%�`ζ��v!pƨ�
�����8�R�S�l�P�_�y�7Ā~Lx*�n��鏲��zp��Y5�_{u�a�H�(F��Q�BUc~��O���q�9T��=��dp'o?#�ϔ}�^I	���#1v�r�?�������@���@�l=�HPK�w�b\bv�������`�N��ҵ���
j�M�W_�?��a�U��yC�%gv|�)'^H�����t�Ɨ&���Ų�� ���C->K���s*I����	f^+���F�$�������7or�H�6��!�I���%�@�|,ڵ(]!�Z��og`�B{��S�!ǿ����O9/ʦ����.{��M���J�C!\�3(?���=�؆	;,���}��WY𵫡�	?�om}6��_�`�{� �ċ\J�7�G�0���b�`7]�q�eM�{���+a^�H^:"t6���JF��
eyȖp��CO�Sg��wvG���S�`��??W��|���޼�Z���8��Mq��1��4�wm;Tg�G�ǥh���¤�|��1�1Y#1�G�� {��}͙�~K��Txf��H)1zN�ќ�^�g2S�e�����x����
h���/�D;"���'���i(!p� f�V�������\Rj�qh�nX���bT8��\�:rz�>����)� �5_����_�CwB�*�Z���k{���߃���t���YW�9bDq��E�`|��P�G�;\oK%y�����R�s��L����z�P�'�q:w%���o����♿���T��t�s6ՙ��s�t����g�n4<H�`/�+�B�ۈ�V�<�x���j�R���r������I�`�7�>H����"��Ņi���]��Ï�p����r��?���^��d4oH���̩��"����}��]�?�S`H�(�u9	F�49�VF�
�j�/Q�M {ۋC�m�G��Ͻ������2:uC!��_��t���,ˇA8{��z�mآnxnA�z?"��<tg&���F��~a�a>��Z��>
>K��K��i�-QP�� ��V��s��I��`��{T�S�`��*��Z�(�C�?Ȓ�&��)��E��2�����Iq&
��_-2_���7�EHp�l���c�M ����g������q^Bwڻ�fg�X_�=y�@ Y+#4�jW� $���c n��H_n�1ۿiV6�^/2�{�a��{������jS��4�b#\{��1�86l��)
!,3�^�^u�aU��sܼR��I}���?����x�>��^z�i8Xgo�L��ʾ�LW��LJ�@L1���w/]O��PB�z���l<��ED8�c�͢�`h �qG��I삶e��!�Q+o�7*�d����.*`'x����g���e�)���#�yu�Ĉ{ ��na]}��?�2t�Q?�~&-�,7���V���6�q2 c�P	����ٌ�J�ﳍ5�D��V �C�O��j7TfNhU�sP��L[�H.�]k��ɛ��W%�w��u"�8�ŰP��Y�p��9�/��X� ��6\#v�(�h��9���V��ĺ�RflFZ�{_&�,öG���!���&�}���q�]���ŗ�n��ʸ�{e�zΩ���r����J������������\��sj9c�Ќ���YV#e�~����w ���O���U'!�<�|(<��R�dc$��܇���}Y�h؋��j��5�w�"�}���FO0Vu�1Q���ܫP�+/���S�=�G�����<�[y�I�����8�q�Wi[i�1�&��,P�ǿ�Sy��pR�J^���E9�O=�zʏd��H䞼���ڀ�gQ�C��2F���I�b�t6�R�6��d�ņ1��>�S�[�rW�/G�F� ���S��/���詃�Y��|�o{R���IWq�:"�~�@���&���E	U��=��D�x�Ӛ��.4�m׿�4��l�oۿd�<9��|�J�<����o۰�FlX�.���಩:Q���Wy���/k�Oܛ�;;�������Y��ݪ^�Օ�Iy��<���b�M�wΒ1J�Q���K0�H�]"d���J�z"q�NɆ:=�ݫ�){�4I�<~�r��x��[���ʻ2�R`��[e>�ng�p�R���X�dK�D�yZeKt9$��K��(�7��n��@M�=8ɗ�3�����P�(�z�7c�ͣ��y���m�㵼1s���B�)��>0�%�?|��ɼc �$'�7�x��O9w22+�Q庐�:TM�T�s�ɇ��]���(����(�1C6��ο�sퟀ�v,�r¨�D��2V�L�2d�kcܫ�W��$��,���I�D��*O�s�l��Ꟶ朾�Տ�Z���2��o�/B���`��'t��E~��Ok�� m������f�R=��M:9xȞ�+9�$�mЯ��%w��q1����Q�C�w�ؑҐ�_��AQ�'���7�s���L�T�z$�k��`����$��!�ժS�T���ж\$�4!��X*����\���&���̻�J@�?Tũ3���]m,Я�>��sqtF2�������Z��%�y��� ����Ѭr.@���m����9����ܔV��:H{�'%Ldy�DR^�n�*KCq��)�!K�M�1�P
>GB���m#��=����@��-�i� ��b�'Ȁ��,��r��]t�m�t�e^�3�����G�����}��B�ǉ����	���Β\�Ȕ	e���~��m�)X�F��;VX���D+��_�kB�k[�͑׀CA�ұ(�o�畂0Iq��~�`
�OP[�}o��[�ǁ���`��hk�z�����0$#�)]32��LyU���U��T�J$эS�l��TL9�d!j���S|��2��R�Fq���y�����紃�;����]�r�0�.��R�R!���3XR, Q���ɐ��"'���� �h�K[ʇ] �|��$C�u���O�:A��m��39��w���Tn���Xx�w%�i퍛-�LB��!�S��|�B+���9���Ƶ�+�Cޫ`�������Vq�õ���ݵ��N�{���n�~
�G�=%��D;M'�H%JP�!�ZB��+K}�/�{+چ�?�	5hOM9�
����ըS@�ZE䄄���M����`Ο�YӶ�fr�LtA.>ݳ�/�/�~s�����O~d>*SF�/װ������B)!%���?�?-����Q6��_�Hq�k��]q��?bɕ(=����+|ps]�;t��-�ĳI�3�g����V�_~�ߟL: �z�;��G�/_Y|�CP"J�ms�-���/θ6K�(��!�OM���8���8�3I��׏�P���EC���H��Z��ŋ/�1G��IzE6Ŀ�[��E�u�{_R�V�� �S:��%���L�u��TJ`F�#GR�0�^���X-1W��|�p��5�H�C��yER��q��<8��XY���O�N&~'j�< \.�O5	�<�a�gd�Y�37j�p�j��xT�7��TT�x�	q�^h��&�GM�k��Q��9%��b*|�fmو ���^6z�F�� b�O-rLRW1'��%����n��~��ȸhY�"ͅl��,�Z.��01r�j��P�7�z�iG���Uz;�v�<	"�?��V���)�'<M�]�'��eg��S�t�%(ㅵ���?�1��_�L	�E��x�-b꣯w���,������<�xls��զ �&.��>>4Q���.W>�lӭ��60��n��7`�}�ay���
�8�B6��愫ٖ�Fx�I?�^�cm��2م�
,�2O��%������΀���<����[ßN��;3�Gi�Y/���8X"�y8<��,�^-�ح{H�M�ƪ���Xحw��\j���Ch�J�����s�<��L���q�:E�[�b���<�k��2�aV�\�<_KxϏ	e�3>�)l	)�ǁ4��PC��d�b��|xb�Q�*m�z�yP��1	I�G���!�1�o�rВ�h��"2�!$Qc����OpX_fFPы��!��T"͹O�\�	��ړ�f�
[��~����Tު�G��We�S�ˌ��� b��Pì2B �q��/�=ci-t�S�$�d�_�/zaL�t�%��?v���i����|	����[̮��En���<�+V)}^}�M3;�&`9�^�(��,'(A��f#�x��e�1�{���;���.Jo�6J�f׶�d���YcQ�C�����o���L���) WS������"0 b��l�z�V�,T/
� ��k���b��O��h�4�ݬ�Z���o���@�(G85�,m .�m�7��W-�Hl�؋�q�x�hq��gBD"���sl�>��@�ql�MF&n��� �Yiȃ�+;og������ȹD)h�^~	ֲ�`���;2��q�y����iF[�<�lB��1�ؠ"dz�Ő�?L24VD*� њ)1z}��WS�l|!	&����cir�<�c�#{�d==y:C����2�S���fL~4����*i���o�g�Wx'��K?�~���7��п9�RKX�+��&�#C��tLz�C,�5����X��F�g<��Z],@q��UQI'�?0�b�tAk��܆)#n���9�oY)-9���}_t[�}b��҇&��hW���c���"�G��4��A��BF K9�~�g�ȁ�%A��w)��\ݘ��m�ã�2�%4���s&7�����,g�U�� ��Ԏ}1���9��\�տ��z���
eG�!���c�7f��zSR���>��Ljj��_�Φ�t2�v!c�hXջ��b;G��:����uB≌X�ʄ�č�RDR������ ,�+�]��S1]�`fD+T\J�WǾ#Q�@�oAw�f?����yNr"2��QQ���j�Aav�,|�m�6b���a��7k)�����V���|`K��.���Oq�I�>�eF��^8��}R���6Bs�^�䙰d��乘&J��X�V�{E��C��&��;�"�.4��㝌�4��]�OX�cU��Y:�ڄ?�DƵ1'h�~5EeRF��