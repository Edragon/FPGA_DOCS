library verilog;
use verilog.vl_types.all;
entity test_counter is
end test_counter;
