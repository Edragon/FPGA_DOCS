��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n���'D�T�t�)�O�o��Jt�A��e�	�zH����E6q.�)_��H�V��~O̕/�H����4<�iģÆ��7�F2zW� ���앲�l�|�'��~r��GUC�p�Yޟ?h��0K-Ŵ{���4,Pd��,�Y$��尞��Ŝ� v�GQ�^�S��9�@��}$����đP���{���/�9Ɓ�@	�(g�֔��X�I2d�o��Ȃ�S�"k�� 4���c��/�z�ꨗ-��5��b���_�:���:~n_������x������g9��ZfF���{�h�5��+���6 ���Ǘ<����8R9GѤ4�3�5�������a�|".#����O�`| �),��-wxp��2�醙V��c���-&L�j�����O4�J6zi�[`!td�	�8���=��IZ��ȴ�������%�V]�IOx���|��9c{�e0֛�����@X��R2��@Ґ}F�Эj��I��Z1��ܸ���"�����C��r$���
;4?έ��O��?��� �
�mg��Cn��;�6j��6�������B�%�]��nz/�Qg�pB�:�"6���Li����k�p�C�z6ki�^�+,mL6j�����Y�.�Ʃ�"Կ���d���u���pB߅����y��i����to��� �����&�a�4$�V�7fP�Q��}'b7|n��P�HM�a[KfQ,��?bA�O�-�U
�KaD^��qI^�����������#���$zAtE�1%������e5VX�4٧�Y����%ɹXN�S��m�3�f+�=^1$LJt�B���ŋ&�NY��|��H�W�mj�Άy?4/��㍺��@�Þ��+\���,�]^�\T�p2S�6���>�"Ü��,�%ڏ=��W�j�^b���4d�����L_�
�u�M��;%Oٓ�لN�|[M����.��4��L�*@Z���|��uF�!�� XP��_�0B�	���.����4ͱ̊`>ԥX!ڱ;��l)�Z)��_JT��qȶf��&U��brbh&z�]ZT�f���~�����Gp7�4wׁ4�ƧМf��)�a��)t?�
kuw!x�ɪ?n�4}�f�Oؾ\����F��$�kD�=3XAw0�ҍ�r��q���
P���1����n\�ٔ�fԉ>_<�޺`�Ӵs�Εb�1�Ĵ���m����oL���{����I��xb�l�����f��pL� ��򘤳Zը 41���(|q�q ��\����ρ`���ND"H�p:��&֔_%Dhe*��Ë'2�Sf�?]�z���=�e()Omf��Nc���s��jCT�� ��[��h��Xe�{����l�-��|���9<ϝY�(���^j����CT�J���(�Տ�0�t�����p��֙�tK� �}����z]ŋ��ܣܛ.I��J��G��oa�=R��J)���,R��# ���ξv�yeL�n�(���H<Xi����r,{x
���i���m��e�F7R�Z�C��6GN�ve����7ɿ^���c�t% �ʶq��Ir��`��n���L�sF���:�:X���&�6	���$(/����F�Z�Ֆ�`���G�� �=��������)�Y��Wbmu����jP�6C��4(��/rM���H�@U?l�Mü:�{q ����۷D�w�HQ��D�\*6P3�4�	@�� ���4�Se��Ƚ��$�8?Ʀ��Rt� �Ҟ����Q�%��L&���7�xȂJ&"/Q����d����oM�*�/��7]���l㣅���j�-�3�&R\A�:������g�����7m����� rY@����#\}tM�/*�%�u�B�k�eEaʅ _mN�A����;�d�rϤly��E�垖4��0ߜֻm�G	��'�ɘp6Ԭ������2ah�m̏�>q��h�=	�U���?�Ͳ�!e��ǇM��W��W��6vdD��Y-��54�9`O��"��ƥ{����_r��1y�;��Uv=v:��#�"�"��h�Ltg�X��1	
a�W&j�n��r�Y�I�,��b��r���Wf���{��W0}F<>��EP�Ƕ��$7�e�É��؊7.��S�毛�/(&R�nl5�T������m"�$�N�Fk��po��(,No�dM\�E�l1�uP�A^3f�&*NW-�&.R=+��b��=�uB��j�"]�\��z�Ð'�|j�0�V��'�|iI/�	�+�]�Pz�1��~uD�������@�a�Ŷ����H����Ҿlr���e,���:��s��5�bJg�y$+��6����fI����ŰW;��:H��=E���1�c�)#�r�ජ),#ڭ���ԫ���ݨ�~	�ز�j芗�w�����C֧@oF��40o��QOB{�+�W	�e�Y��`.Uo>����F��/@�_T���t"|2��2�Q��vᜇ� ���e���h�gf:�><��oQ��`\����o�o��r��#��ޖ�)�x:*z%�%��'�շ�c�g�=�V����I*�9�%ϖw���#��Z������E�	�]�m>M�����c�\�{p��ݩ��"����u��}v֢�����7r����N���Y�1��hw���7�����(d�H*sْeLh�@�:��ă��5k��2����#x0���;�ZZJ��f���|����cf$�I���~�(�X��N�.��4�{S��$���̋�Z������Po0�����"vn0�\�M�a���"��z��v�X m�[��ʊ���Ji޵��0(�}��%1�b�2�m�����J�q���<�v��m���h����S�i�2��X�CLN�i�|\@U ��@Ω��I�H�����I��S;aA�Zm8貤�5�m �ܧC�X��CK��;G�eKD��CHY(��\�(���ޑ�wX�	s{=�rg�!�6{'m�*����},,�{�ꆽ���{͆Ô���!a%�pq����C�����R��L�'.��1r�7%��Nb��:�x�fW�B���隅�~��a�D�y�']���wd���^��~�2=u���=���	CV�V����D��KQ��|���^%ڡCU�K"��]�ʗ�������F�G�H�y	j�Jw�q�@�����{�\���a��|�׺綹��cN	̓�ݤ���l�(���ԙ���Ƥ�-�Xs�o=G]5�(�ﭛ�j��H�����T��Nm�Ѕ�z�����A�4 �Wzn&^�pFƽy�8�^US_�Hz���L��N�2�{�ɦ?#Ʀ�fo ���&�B}�Bn�*�����|	���7�d���ࡴ�(��v:��Ѵ@��NF޿�#���ǻ���=�Y���7m��JkP)�����ݱ�H/)��d �t!�"lw$�Ѯ��+�������<�߻I"pw0|�ce�a K�ߗ�c������%��:W���H�0��D&$Z��x�	\���yJ�P��[M�\�彥ƠǮM$�5tS��Z��OA..o���H�Þ��Y��Em��s��k#+��#���:�g^9�!Ȭ��
��
�-�nf9�b�s����l��8���}}���fr������������>yL'�K�ƽk��d2i���6,�q�Y�)q��X�ra.�HR�'hb44�~���/>қ�6��zhn&Z�6k���p��n�͍&���B��/����=~�<m���x�u�E(���~�ͫ��W�vTGB����&���2ˀ�=�DM�feOd��&��Aٛ0Ƿ���RQg�D�W?������j�4��*��z���ٙ������4��*���	G��^�z�RN0���#�C]�*_s�Sm���G��2Xa��?��5��sL9�������x������D7T_���ߞf�'�p}LC��H�J}�x���C����!z`P<R&�?���|8t3ԀJֈ�b��w�S(��He
y�瑳6�P�����p��^v��܆��$K	��ө�`�A��n�����/-��A�h1�C4�ot1q�5v*;����iJSs�D�-��H9��(Ҷϟ�+�m;����EY�es8���2B9��n��e=�M�ݲ�T�9 V���|.	�>�a�oSo|��۱�Q�Sb)*^\3�����k��w�P6mۆ�1l��̪� [�J�J��:5�i��j�)ʪq~�J"/%�[R=ّo��eo��YB�{��3(�	 b�/��P���O.ӊ{X���p�-{���L�����֮����[����I԰��� $ڸ�T�dQ8��֑	�8�r�Lj,�d(��ELc���`b��c��C�8[m��1t�xP�I��e@}�9��7��A_��u� �m����&�'����HY��c��+���iܢ�����5�T���2�El��>/<z����|�ɟ?�)fk��ʝu��B��9;�h$���;�((�;�-�W��ԤU\Xr�����W����M�+(	b���G�Z����>�����	�� 0 ۏ�ֲ����5ݳ穻�)�{,������ă�&
ٚ��'�Ec$��P�%�r�����L ±�sw�Xd<Q؝Z��~Y��S�KD�3���������%H2dGB�#�
6�ʰ�C���N7>xB(��ԉKL�y���Z�c?`��u����&��0VT�M����x�?�9�&X�s:U��Axiށ�nq��M�ģ��@h�̘��DL�K}�$A��*IA�z��e� JP	�J�H�M�
�F(���Mz/��Ym���IʊaK�	hNu� /3���>">2zƊ}L�:�(��c�����B^T-@M��gCjr��d{nw��9f��j���#T��	&GI�,�M`� c���e��޸ɽ�t�MsY�>��?x�m b���u�hy�,��<�h�ȡ��=�T.�G�;r(�EA���m��N�\x�c%��Y����M�o�� h��L�P|�7��E�;���.����/)�j%��̅&�da�1�=�r�
���
ԋN�����oG�{��i'��fݲ�(��q.|��^��x,�v�f�ҞX����s��K\����*���o`JS�\�g����r��:��y���0z�ĕ�� �>�2�2���@~��m��e�A�v������5�G]@�o�)�G�B�U+�n��TΰMuIX}:�~>�쏔d�k����N���tJ5���?��1فܲMN
Lf�Jy��J��C������C�OE����g�1�u7Cv���6lj �7�� ;��[;��^��^#��<w����Q��������U�=p��@�~X�}}8��Ow 6�4d?���z��ҟ/w�l��^FT7�u3,	�H�n�yM!-�ĺݘ",S��'�Ps�@,G�����}��X�it;��/U"|{��|#�&�j���S=����w�|��BY�K��,0nPG:r̟��2��8[)L|��I?��d/���%H?&9�u�L��@IS�����$����f����,d�5<�
|p>��uډw��:&�C�z7\<.E���:�f��M�L�~��Ϙ"6$T��|���|xհ�^o:{Å[.H�r��ϔώEt@�V���n�n�㣁��z򟜥f=��\u�c���w�t�{�Ǽ�	�W>�!�l����w���[�-�.�fOr�>�ƸM?8�הV$�Z!��9�X���wN��q���ZN^��8����o=�3�3�V	��H;VyU�� �V0m1��q�j]&�5U1!�����`l(�Q�� ����r�bۄ�5�q�oK�F�&uM�«�J�Zϕ)�-̚���ϊ>�h�� �iD�'�v7�S��|�d7������dв�0�{_5;w�RX;\+�w�.W�G^5
�ib���"w�������<�g̫x�8��q��W���'ʑf�v�dy�x����e)���'�[�8���h�O�� hO�u��7F�}��6@rs'`I���T�h��g���s��C��'���q�*����C��[��А�J�+�d��j�Jl����Md:  EQ2��/�������#�N$���=�J0f�Ԫ�,V?�(v���K�E�E�K�d�����_�G���C�r��
��A/� '���7�쮒-�;%9tY~u
�l=�M���%�1���'qЋ.���P�ܚ�Ǘ���5��� ��Ӹ�8� J�=x�<��7��q:x�� 0�qDdI�p��FJ�]U�� �'�R��N��S�_����T�~3�shf�֗N����ί~��+ߗH�~�Ye�}�1��V
�6	�tȸ�U3��7S%����~�a) f���Ց\u��+��D��T�Z��;L%fq�C�.�c������s���Z|��}&e�T�rg�;��()-��ZQƚ������e�~fp�f�6�Y�YB.Y#��8)�A7����͠�nw�[�(��@���k���d�a2#D�)VR%����&�W�*Us���U����3�t} n���bG�
� G������;��R��8o�]�UEi���@�Ɇbםw��%������(��_�Wo7�����f����:�HX���������֭g5�!���(��r:~�R�N
 ��T$h�Њ4ay[2���*�8�T]<��+G5�3�������>�%�_�Y�][۳�&�� d�]����N��=�.�l�)��u��v�3�c�8��*"[~&�亞����G�%ύ>�^�	�m|����/��ϙ��!�[z�*wN���C�j��@?��K���~̆��]L Z��H6Cl�󵔬{ׯS)�y�C�k�`W�>Ku��
Xa���{�HP��[+�@�٘��e�^ٗ�7�����*�ˌd=kEYĳ�h )�_�?�g�mA�hhb?�RZ�'��DZB%�R�:Y��]��]9	���ط�3�M��Ņ���EV+v��׻����T��׺��Y�68�r�k�
4o�d��J�G�B��l�ߜ~��_ C�f4�c�[=I�EBn�����rK�38K$W�����KP#E�Wd[��"^��~%D�X�I�J��u�3���-���14C�-�jZ�s���p��l����!�QK�(����xၯ}s�:�Y�i�d˘�ue��E<�)���9�3􁃰���,�Yl0�	�_�d9�V��9[!0���P�����NoWV}���3S,�����[�\�wC�`��ڄ㊈Y�B��D����D-��]�����b#��h��}�0M����s͒��UZ<fd,����G�s�]˯_R����Z�K��K��V�݀	k��t,R�S?�B���R���[�т0J��w�d�wh�<}p�Mw9��L�V�R=�}�����d��ͭb�����/�XtE%�D�w\�� �����P���]�^4I����l״���G�����&y*�[L̰<��v�aZe�ǭ-ȭ�^��U�/��'bG��� nNJ�sJr�j<h�ve�q]=]ಀ�{R1��䀪G[�k	%1r����vB{�5� �謾��Ў�0�c�3v-#ۀ�ܮ�|� �ȫ�2�;	�`"��~�oF2i8O�M`���i�	2(b�UO�J'X'���M�61\Y�U��a�Zи��Z��3z~2l�=ɹ�D��-[]C]�Q����T�4��$�r���Rv� �@ΏP������+�4T���پ�{K�e7��~����[�xh���|��w�C�������c�l=��G##����)�lt_��Y���o���Jk��S�#�V�'E�"I�a�)h��O@�~���:[	䜌
\&aE�R���_��䋖U^���m~�T;���o+��GT�t� �t�
O�{����􏶣Rf���ڔ�;�T��v�T�N����ѿ�ꮒ昨��!��� �DH	��	a�G����VˇςY���5��qB� Z2Q�^ɓ��a4���f�c�k%�U��7u��^��'����^six����=����4�4�ř彚�:�X
�=�!s�F�����|5s��nB�"5Q*H��آ�}	t ,� *L��C��:���qR��� �O}���g�^?�:� ȹQJ�%�Q�K-�1.�)^�!����1���,�`�d�zC¸E�:^�b�7�Q���V�"x0,W�$q�'=�P��!$�A�Fz_���X$F�m�d���� ���B8,�5գe�5�i|��<X���:�lPY�U�>��Oz�g���������/��ݵ�	bڜGH��Xs'�ſ�>����p�Ɲ��7��L�D;�#�w�L�q��{f'��Ǉnco�i<��M�P�8��x���13���P��6>vU����ހ�2c1���{� ?�GY6`h>�&N�E�'��/�9�G⨾v�N&��f6C���|��z_4" ��W�c�I��|?~ࠖG0�5�#����GXZ��X�T�����a��K؞B����M�0�����R����A=J0�/���f
��h�4�܌r�K���|g��f��<���*%�z�2&�$�0�km�|������K��B2��1e?�<&1PK��i%�3�=v�{u��Y6~;)�)	��l����%16i`�y�Sk�����m������:��[Z�W�����X4�@̟�ȨE��@Z"f˒R�x4���@�	�E�%�����N*���&Q�����v���]�[�IX�����oU���C�]���zyq��Xo�,��T%v��|��<EE"{G�"1���%F|�P:���c9i|!a�i����a�Ђ�����!nI���t2;>��*Y������A3,?�`L�w+$����7�(қ�Պ�������,�H�Q�*0�1@���xǠ�,sp�P1��F���xO7��K�o��~�[i-:�[��}h�fJ��a��z5[Ö�`��[�
(�܂��m�!b����Tzk��i�o�y�،����i�4(𿕆�oh�A�/��:��X#>�@)1���:�1�J?E���*dm��J��ؓ�25V�Sݤ����[Io�#G�%Zغ�Ѫ��}ө��ڴ�&�����W{n�mG�~XΏ�H����{���}�0���v4���ɰ�����X�nM!��ຩH:��Zy����� �<��&Of�L��s��[����V*�/�P�W-���W��� �V�R����B��-�:a5��p����G���R2�jJQ7,�d�B�	�ϥ���-u⣦�KX3�ꈺK��&4]�#w��%4�p�Q�sW>�C)��Ub8?v^��9}���Ag驮~�]�I�٭�%X�%l�QMĉS"�0"K�n�ytS�9�4�+������[q��4-�8�4���:B��8B�Fѻ�u-�zז��x/0�`�U�wO>�fG��iq��"�Gt�P�4�c/�0����4����sE�PR9;?i`AG�s�%qmx�^�ԦQ�i˼hR��VX��{��_�7�5�G���c��ð��._KՊ�7:��V���M�kON�����\HJ��@�B�DE��e��*�&��S�A`�we�3�%j�e�բ��h�i�Tf@��2����SAއ�P_"�1%�"�m�Ǟ"�l`I�9���	�٧^G�6��}�V��]�|xIρ�H/qs����c_��EוI��:���Dl
	�d����ʜ�D�D�_�h~���Q�84)}c�g9PzG.�)b�/�3�L8����Ɇ�ʅ�
�-�?���	�j÷�J�u�6����!vx�Pp��"�а�]R;��dQh� ���~��㮸��Q��%$�0·�}�y5�.*V5;@�� y��k�=��ɪ��8ߏ�^��0��̷��;+	��Em[��r}��#�]��Z&��_YDHJ���|�b��gC��z���&��N���@���݈]-a�Y�bh�O�$����EqK����w�i咻�-�;
�ϷXL�� [B��ȧ��f�k߉�xw��
;>�#�e��m3��7�~6W��~���<���Uyg�č�nY�����2����(��lԹ���Ł��:#�GQSV3����U��:�#����P��y�@�2\�|w �+��o�N(�"�:���ql��׷/�����S_�#�Jk)v��-�O��3�����eޮ]Wy����v˨�r��/ɠ�K�����h=��P�'���F�3�K�r5���D"d@'2�b�m1�eqϔ�&bT�a�E�����Td.J2`�7ݨ3_ժF_��F�.��(Yû��:`��^�$���D�y��s�-�v���-���.Wf����<M��5  �;�7W,%����B�l��[�9���p� ���΄ص���A���]�9P��֊0�3����[�q��$F�zbߖ��)���Lp�#m�|�8��SUt�Lk�z���wG���o$Cva�W42�g�����D�61����&t��n|z��҈��T@�A��$�����9�t�'Jk��N����c�\+�"0�B�ٛI*�\���@,Ϣ,��4?�8A��6��w�A��Z����fM����j��KNC��.�L��ѓxF͈u9�X�����#6����۠^����Om���@�Q�ݬ���o���T��!���X�'U�����B��Ri$i��k�X��_d�W%�3�Yo!��&I5����~p��8S��Y�>��b�&���-a[�hhU��PG;�Ԩ�F�(N�R{����27_�B�h�l �H)6�ĵ������K��=��7a#��Z�E/�`%�� 4l�b.�S3�i�ڊ�hs�L�6�YtY?�V%viݦ��(����y�$�@r��H~��$�@1f��V�Ke�c�K�{�$�F٢�Č�>&bm�� ;]J롮��_j����� ��=�ڲ^�B�"dɮ��f��'�ᐚo���c�6Z=I�������8�M>��#/����)2��d_�չ����R�VH0�pG�`��ߡ�&�wa�<^�le����_!�=jA�� �,�-A݊�Mt��c����i@���R�_Z���q�U>D8�	"�.�06�f!Ertr	N��
�_���N�<>1�����!�JU?^�Yk�>�;m����<1W�ux��T��y3��4y�����Ť���-�z��TJv'�T�ӄ]�LwE��8`����~��Ձq'���SP3hq*����N���Vz,?m��7P��+s����SIS}�m�$��v�	���e���ֱ;=I�
�r��Zt��^9��Mw�2��b̡;�&g<�Z��7:��BE?o.����89��7T/���h-�.gh���F2�b��9b��\9I�l.z��˲��N�W�4}�
Y|ſ�ߐ�W�И��K&��b��q5穵�_�if�by�B�7�8ʯ�;P�.��ڣ���NE�����	�A�2��H���g�����߇a���UYFL�K��Q�?7��{W���E�ͬ�<yC�;����1tNH�~5$B����GYA�6��MqL^�΋\ųnE�
$i���[FBڢ�Ih?�'�<;{��S�e��9�
&taF��;�MK�/�-j��K_���3�sR�x���z[�&ut�`T����,cq(��k;U/���T�[Nr5��R+_���T��f\�;��N�cB��?�����M.Np�����9�/�U����Ĕ#�S}�������1��
�]@y�qa���i�c�c�����^�}�H�4+[��M���6($��?�Z���U<ͯºl������48r�{:�.�F�t�o�S�劊�ۓ#���s]���BN��2��hVQ5cyq��t˭�`.�"̰� ����pz..6�7�J�����k�妵_W��Jb	��^~@;h&�T�Uļ�⦹$�5|�&k�S�O�H~� i��}���\N'��F0	˽EmR�����O0�1� d�ar+��-��Mo f��^��ʮ��sS�M.�v����	}H�{
/8���+��2�xCjw:����8̰��G�t� E��?��6��1���x:�b���fʡ/)sq{�wN���z���1s�%�m�i���Bq�������f��"���E(�Y���`_�r����p]ۊ|��x�.X�ު9�z	����F�
Q<�M��.�^۲�����@�y#x;g%���,P��#��q�"wP#s/�Xlq����њ�2e�$�1��r+��KR�8,��6݊�������ذ��!Q�R�62�6�s/�Fpk%��"��R��!ɂ��"�,��V�����6�+�x��Xg?I2�n���nq�tݻ.�V�!��zɍ�aX�V� ��z��S�[6�?�^3"����oj�h�sX#�c:��L������2�a�YN�O�5�H���ɦy<���[i�Gl��e�C�3��^�S\^�������.t�GR����	'7+������p�v#Z��Z{���L��[� ^���d�~�홱Q{��@��ɇ�;x�:ÐR��G>��ò�ìR\_2�yn=]ȓ�V"����{7�,g�T�=@�'j��.9�@9�q{�M��_�Cr�]rZE�Zn	�T��u��S�x��Ι�H���o�y��@Tu��Fw�ljP+�f��fS��ƌ=H��n���3oŗK��nz� +�{�X{��jy�̇x2	��=�G�h ��-�0��Q���O1E�*œ�釲5Z�Y��'Re$0V��G�.T���3H��i��pECQ?�gK������
0�=��i7�ɤ�� 9�
*�]4� 4��Yr�U�;�'pǁ=J�w��5m)Pٮ���U�� ��i����P�_(n�x[��������lמ}�i�т4N�UW?���VrX�B�v�6�z�"�W�n�'�V��rP��ԉ�L�@-?�0��lsʏ�ä���"�~6��~3�G2�rTJ������,+��1z"�?Q'�~l�O���
�����+I'P��v�Ģ#�z��y��k�d5,�'b+20�+��T%6)�wU��8yD�ge@I�Z�jZ~ �sñG�}g2�Vs�=�΂����I�|c�4`8��=�Z���HH�� Z��|Ӓ����<r/������Ǡ���1y�v��M]� �}|q"�� ��J^Hgi5u��D��܎����.��P�o(Mc��eoa,��V��si�(�9��К�,�*6��g�����"�^
J���;�zS�MW	�1���ʖ����!�G|�������ǧ���f��އ�~�x2�Ķio�l�M1����˦k0u&(���j.TG8y J6�q{�8"C#�,�[��HSe�n��8^�Vfj��6B��8΅����z �}���� A2���:�WT09��#{2�	}h
2:�ql�͆���}���^��i��+o	�\*{��`�<l�n5�.��X�e�5ˣ恗�P���%��n�E�e�})Lō��޼�@��
��z�<�Qn,;c�	�o���	d���0Y~�!IO��5��2d�$�uH;ȕ�>⿒�ԡ��܊�O󚕒�s�k%,َ5Is����%��U�����4@��(Zf˽��j��A2�>�w���{ e���7�C7�1rY�c��D����?G$�h�#��..;<ޢ��p����Ok���_R�vr���aP�Q�5Il~qB�E���m�"r�A��כ��S��fW]�uj9Ƴ­FՓ��E�7��%�+��d��xYw��h�\d����R�֯ϰ� W<μ�X\�p��bb�O� �%�(�X���A�[倒�kޅ����ԭq�%�i�@0p�9�,��[×�����_�d]�$5���J}�#T]��$� ��;j4�K�����Y�	|�������Ra��X �mu�7 ΉQ�l�^��N�Au����1^!~��j���F�|��t]�׬�0^�ܸ�k�#S�Yf���j�~���T
��O����R]�ɚ�8�fj���J[-�����X��>�Qd�E�����d�]���=J|ى���荧;*��g)�>fJ�}�ۿOj��HO<,)>7Xs*���m�c0��Y>�M����|
���^���7�T�*��du�������#��a�!Z���`����� ��B��.s�c�����l���/�o\,q�U�b����|���F��5�"��V��)�41�7)յ�q}[T�Z#��
���A���J�H�Ar::q:g�P�V���S��gec<J{��#i���C�bB��Ȯ��4�U�yX�m ��t7����G)������U_I�1��O�u=5b�1xb��(�o�y�=����*W��(jӘ�-د0n� O�v�W���#Ņ\g+�*!��[:�
>��H���V�E.%{l[�0���\�ВKpM�\�8�fh��^��Y}��u��2z�-�-�&.��{H����OT<Z�͜��.av�۝Bd��)���xM9i�|e̯�"��N��4�z��(aX��0P�<Kdy��	4Gq��8_�*u3�ܓ)��M����g�j��k�/��J5%�e���@a�L���u����m�(<��|�����u��h�S^@c��Ө�
��}�E�\f	�?�=C�.�����{�0S��w% ��0�\0hz�ft<��+�Z7A��0�O -�����S�\�&��zGLPi���6g��v�JEf��)?!g�Y����t���������GgI�&��{�����E�3�oɨܨ�[4:b�Z��?��ɬ������IQ�|���V	a�+>�]��!�(w�W#��C*�$���r�!3��l�t'3-q����Źo9�|���S�`U��Jz�#L��UuyȲOH��ˊ�S�]@�'�T�o��]t�����A#іy�1�XI�aT�	 �<���ZU�ڄ��j�8�H�B�(�է������^��^�2�2����c���_����ؤx/d�r*�k����?��c���z���)�L\�%������!68�m�cl09�*C�8�.@{{��现^�e�>���Ǟ+�,�y���b�j3������ R�gJAj�KG�I.\�0`9���̸��(>�)�\It~
�.i�aj����Fk.D�&Ɉ	W{C������m�`/6;=`c�p=fM8�
Y���C�_
��H�>��1s�/���w�Zi�E�/S�>��)�Ѓ��:�"�}P������$l���Ge�Bg%���ȭ4K����z\���r�$@��w�bnR �� �0�w���N5$���Ңz��U���篝h�oم���U�{Q�G�BÎ��D���-��'�g1�o�t�����H�p!��5����[��/T��,��8�xbu]u8�-�,�.�7|������?tD��簴!W7x��)��$m�#�����?&�:Xʙ�R���.��- 0k5mz7&T+ :�[w��,�Y�`����Ź��dx�$;+�������e	]U>9)1u/�l����Ѥḟ��6�w�p(�N�~�9��g�MJ�x)��"��!­�����T�l��I��.�@�W2i;
oŷ�F������`øu�KKN	�i�߰I�>��UNj���b��Fr�@P�u��1��E����+5��d4��/��di��t;Y�˖���%t>����Fa�:�h_[�J1�����^�ͳ92�9����[�;���~��5f��+ �h�8�IVq��Fs�$=���a9��Пo_�$:˳f���Q����L�B� �~�y�$l���q�r��1�i�t��F�y���2or�߆К>nFNP$��w9�7��Nc�#GZ?Y��p�i�q]��H�,V���n��FD��ڃhdN"><%�LA$������P���j�Ŗ���E����}&�̗�[�/�B#�8��SX����<�RkxW�  ����Yh�-��L��_}����+�(�1׻ޣ�z���Y�?O�k��u�2E��4�QH����o����$������ ���,b�Vކ,t��T�?6\OGHՒI�g�����K��]�ժ1m�r�?���;6{�R}(��Pz�!K���xB����J���D�~�C /l6��B��=�O����ͼ{��׆5�dՉN�����W
Ȃ���+�XA08:��r�bpF!�Gn�,�,v�N�B�,��۬�Q�F��oO�δ庆�[8�b���q�N��h^�$X	#'����y]e��jk���C���#��Xb������l���5�t2�����4Z�,rʤ��5��#�-a��.�����Ds��dפ���2<C���a�3\�E��0_��BG��$��M�2���(�j/�@|�- ��J-��a�ǉ�� <$����kl|����'�?؀�I�ڃ�����G�h4����!a
�>-a�J�V$Z}WU�sZ+I$��;�s�cI���

G˪��d�p4���gD��.�0�(��BP����N�"�u�,�)� %ۘ�/XW͐}Jw!����j�G�F�z9�RT�sTH����=�yM���택-ToU�!9Y����
��6,|'��2CܢW����)�������kk>�U�D���H�e�w��=����p�b������8PNw��)�!"Op�;�:�e�tl�S�1��� �nK�<60��9�d-� R[$ra"I�L������d�I��� L��{6GC6�,e�՝����4�0�>��`�f��F�?=)�8\��C �m���$@\k�������;���O�QBg��w���<m���}�~����np�g<�]�Sa@�{�g�Z�T�<���Mޙ�*5��Y� 15V�΄R��ϩ��\�	���>��"�&k�I{�5vq�)7�8W����M�8P�=��@��������w���Si���a�ax�iP��k��L�Q�����y�L��w!N\�^P�&�� >i�ڙ	-��d5됎$�Id��#z�:Rp_���BV���?���.0o�Q�WHs����|�����0x��cK,b�0ԏ��;X���V���+���'��F���V��H�=㠅GL{G��G��,�>}�����}
�h~�|�VP~�q푣� ����~1I�y�a y����ơ��6;�'s�y��K55?rJel���v�,V�jKAi���
�c�h�@���Er��Os�ol�\-�=;wBXw5y���
����?��Y��g�O��dc���+�3����MK3��Ƒ�������X�±��'�S=V� F������_��w��p�g�Q�Xl����Ū���gh>��lv�H^��uX�WM%5?di��� ���X����d�&#�G�
�f=�@�x�u�`��-�.��V�?)^"	7�����_��Ifd�]秺�A��T k�R�.e���??;=][��{�eK,����W�&؛�v(�ƌ�Ο��ׅ���g�Bi�S�׆��S���T�IX9W8{mNoűF|��t�t7T��ک�C��T55q�(��</1��r!3���4���l�#-��O�?j��ʐ�Y�7�Su1|���~�N�*"E�6m�g��1G�ūK�U���8�[�i�fBg����S��λJ'e����/��ָ]��x�#�Cf�&'�!���#>����F��c��:��A��v��q�v�����ky�MĂ�<PҨ=V�Q��
3�pZ���)�&c��=b�,M�Rp*���BEnA@�#Q"��R���}Gu+KG����g}> �	��S���Q�U�xt3��*B��o5�<r�Dc�pLz	��PtQO:�����/�86��]^}�(��)���#W���4��XC��}+�%��m�)�J^n�1B�j,��9nQ�(�{�H�a�i�a�U��9o���D��?"��t~����d4.���k<|�u*��t��j�o䥒�%�*��C�����[���O�Al��=�GY�^F�Nx�^f��y���s��l��F�g�8��9���K�Z����>�[W�>E�hz7M0֫�eߘ�Xm40�+��AEm��[��/�u�/ë�̵lk�����vE��ru+���n�����L�����لh��R�hH"K��{�K�����Ց���WZ�
3y�o<Ҙr�D?]uvy���"�Ubj:��1��f��S��f#�l�C�W|�q(�C���*B#��~��C�
�v5'Cx7��aQ[o����hAs�x`X�g�\����yN"X��C1MND�����?���5֯	��F�\�����x�IAGW��y�ݓn�X��w�����{���j�������WE�> �tr��RyHkO�J�W��`��\3̐ ��p����>�����&G��X[<��_�T|�q����R3-:7�,���/��Y�}w�����lz��-�B����dl5G;R=8����E��P���ztlu.\��}ze7a�5���h�S�Y+ F�]�\�r�WG�)X�=��3���Tc@��Ώ8��#��S^<�HC�p�U.m�����$�j�g����g���fbv�X��/�oɩѷ�0�l׏�����%�-�����C�g�#/�b�ޮ�KG	/l�izë wz%S����x0{�94 x{Z�1�bW��:�u>�pֹSR4h�B�������-M2��7�4��[,s�K�J�e��}V��*oO�-ӽ�'��?~�L ����.�.�&I@c����e̼�9JvW�, �C+(Y����N
`P�83�oK"�Th�)�X�F&�������5�����	' &���Q�`/":�8�
D�8��|�`�,�h%�	�Z���Y���~�*�<e��aј+�d�0�;�(��1�~g�s�I`yrMT�Dw�z�%��
S'R��=����L �3�dk\8�h�z����Ñ��*�݀�<�����y�3fc[��������b��"E�e� �b$�]�lB
��c<b�e���r��q��nc�H�Em�e2f�$�vX������R�n&�m�	�`����W��.�9����?̀\4l���2�����}.)v�s��%3�>Ey�]�0�@l<~ ~��︪�TuI�"[��
�����꧖�m�ҍ��n�t
Y7�v^ax�ϗ�B,���nQ��mܶ�wz�(o�N�1����c�yT����PK]
[����RjO�W�8� �d��{�H�j}����3'.�M��-ǙZ�mu��EH-j)#|��i��Y4����An(^��:n��	���b_�͜4�J����`�)��=� 3� ��~*��@	S�m�:']ҞO>)��;�M�?��Q�*�L#O,z�\p	MU��A9���9n��)�ϖ�1��#�7�]B��+��WR��\����d1�y;�S/�EN�?��⠡AdE
6\u>���(�q"s���
w̮�II+��*�CR˙<zV@ /$��[����`&~�N��=pD�e(���/S��Y��Si�Uŕ��di3-%=���hz��3:jOQkļ�+��SG"�d-�|kN��&��:����������XKI���[4oƞ 22���lT���������,B٢�!��w2���Y���sZo�dc��+,�+߳��.G���Q=��q+i�
&�ĆrU��''KP�$��=�Cꖓ!$� �x�8Ѧ_��FsOɄ]	��ۂ�KF�W�j�{��e�\e�^z�O-�I�OB gD��C*�M�q:A����/�.C���n�ܨӓi�>�Y�#.^��`¾�V�Y^l	���lC�(F��O��r�q��ه6D��������0x�׹I���(n�-�ɨ��E��
�|��9ZՊy�x�׸�83�ʛ�������<��|�)��b�	��;]�D�F���q�os/��f� ǦW�Aڊjs%}��\�.��P^a^s�C�w�!*W�����+��9F��,s�b����#��6��p.�޼]=�m.0@��R�����kRo[�1���s�%��t�Un#�(;��8������4���U7M�K�s.��̦S"���d{c,��ǳ�}B��N�=�D�F�B���R$��7�hȀ|���p�?7��������5����v�WZ�)�A�xx�j:]� ?o5[���p(�=t%�A����C�{���8v	����yPK�!?4Pc�T��9�ټ&P2x���x�xEk�� ;�uy��+<�ϡ���wR��Z��=No�+÷LV�����ƞ]s�u�	F7��/�ZB��\M��c����_����#t��ƺ'��S�)y��(*#]8J\cMH٢:Ì{�)�7��U]�#���#f�jt�ym�h���$~���b���g�^^/������A�Z����xJ�)U��
�-�^���W���������<�NR��m �n�Ǘ	��h�1J!��z|,ee���\W������A]�PZ��0O����_�rF}�q�;;$��',�_� ���%v;�s��j5A�9G�7�S�D�t v��s��NZ��u`�s3���md�����  2m_7L��o��&=���LM
c(��&���n�Я$�@�̓�Q~u�jj;��*��x#l3�bEJ<�4��F	²�������c�H�d��?��p�q�c�4�@�L�`�`ss&pi-�^u��|51�@�p�"4�B�x��G#-�F�.;�$޲��-Z��Zke�87��v���b	Ĩ�����Q�N }>����֐���X���L]^a)����J_�w���VR�x�S�.�r1}ք=<����(��$/�I���X\�&�g��W�k�)C���͜/�z׷��VtWc�'����qF�ʊ5G��яa3��J$*�Ǝ�eR����a�!a2R�0��/�
��O*|�51�?�k��q���L������D#�����(d��Q�|����w���>���a��T+;]�iW[G���lɡ��_��,��b`�`p6�@�E�7�㲡5l��p�5Hz��'q\k���x��95ИЖ`1��/���{�)����Ժ�>��;BURs��ξӛ�S
�>Ǡ�@l���h�+���I�0���{�*�Wn6+��o���5���N��B�q0��A�2S(G%aV�W���h�P���)�iW�� �M��7�)�I���_�//pJBF|��o&��0΃H�ED1�	JT��j���~S:ۏ��G3d �`1d�\��g��&�*e��3�Џ����t�#(
�?4�p'<;�Eh�r<�����j�b�_?��r���L�0O�aի/��)�����仹�7P��!ǝ¡տ�~5{�����0��Q}=�"���K�I��u��}&����M-V�O�#��n���@o��+0nPՓ>F�:������WYkr�!h�Ä��#��cز��.am��E�`�~�1�&����A�����L^l�uN;
H^ݣ߄��c�Z�4��I`?*Y�e�+_�Q#]�!��t�ӵ�;Z�ÏO�ׇ��V��>6��Ɇ���jR�=~�hp�rq�XH:-G!�ql�/�\�{��a������0`�`���������*���t�A�NW���E�T��EF��4ڬ ���*$�H?�������j��]t�Rϟ�f�	㮴�����@z�/Y,���?��E��[�D���F��6�"��ޥ��ڀZ2h�'W_,�
���ID���>�����_U��W�s�O�x�����&El��`jS@s�ӭ����9#����s;�ڳ�{U�`�R:��B�����=�h9!������	h��s�0�^���)m�	��0=V&&��6�B����0c����_�,�RG��Ffkm�-�zo��@Y�3~�p�.y�e>��^��œ���߃F�����$�,����4��a3��Z�Ǉp�X����ћ�_:ˊ5�U%~�x��ɛ2AӒ��j"xѱ״�m�/�O`i���r��({SAm��m�� (ӆoV���'I&o��E��cxm��X���(����k��HEu8���ߌ�p%���y�¢ż�o����䶭�N�%ѽ62&��fP����G�����xy�����ΌI�.2��n n7vԊ!E�	��<$&�曞��G��\G>��'�,���=��p���_��1?He����	�i� o�CX�*s$�.�;"Fؙ�r<;��
�4Ǒ���~���nJ�Uz}ѭ ���)\;8����/�GP�#J#�(d	Fm���pO�^%0~oBv��W.W���  V�җ�9&�=����q��tXYrt�̉#��,*ݮ�Z�-�a���0g<�M�3[�R[���
�L!�mb<2�_��Üj�4���q�.U�=���&+$~�<����������� O�$�ObSV���[����a�%����ܓ��~�O���֍�����U�*�̝P�v���6l����>�R�I��CGUʬ�ˬ!Iڒ�����
ū �>��Ք������$�d�#���UBC��G,�lrc5��5N-���t
k�gEw
�sZ�����Ͻ�����=0�V�գ��m��������3�)���9�����BU�Q��55$�,r�=�r����{��z�?^�7;Н�E���y@˟�����Q����~W�B�7�麕����w�v�����/nI�I�&���G��M�5��� �*@-n"�l�"J�]CÇ9�!a��֝���mQ�-������	gw�W����2���
6^tk�ֈ����,l_���_�\��ƙـ����W�a���K�/&�}�e���%�6��bP'��5�"!�+{�,��i�l�)s�F���'�Tܝ��ބRJ^�.#wq��jp�<���1E�2��+x�/N�z�MMN�n�W#��ks �%�oI�$�ބ\4
��l��*����!��;�#�!p`��5,��_(��^��=��7��'Zrs�� :��_6lL�;�y0=4G>��w]Q�G��� ��S)�xZ�r�9o�J)�J_#����L�ņ5�s��#P��o�mn磰�K��(�qb6~�^��A��R�W�%����bt<h/E����l��Y�C����zs۠�_�(,���]ɆB�y�n��W�溸��R�{��s^��jwq5�䙯�?G!�_��M�`��Q&4S��.u�쀽qmI	�I v�y Cs;��ys���8���m���r	� �Ǯ�����j �6��*�Ѻd���{D�\�!
5R��Z*�J� �����~Kq/�eE>jY �5�vB�5�+F҃���GZ`�d��ɢ�d������.��	q��g{ѵq��,w�Z䄅�S�M׵���iD��ub�re����ǰ��u�2���쿺cі��*$�����#�:ʄB�Wƣ�>-���5,!��i��1�� xd,�5*��p���-�ST��~Ȇֲ��u���k��"I�}&��#����n�#��݊��k��߷2���d�@��?��2�VP .����Js�UL���)}y
.ڙF��
X��v�z�]T�\�-��w���b������}�'v��)u����%�+�jW�o��Ss���k� �4����-Lp�90�����e�q�Ct���,��)h����q(u,q��/q~`.����j�
\ُǷĿ&-�{�����1A:d����S؊&�7*��c���������ձ�7I��eq��_cjK�dj)��%#~I4��8&	R��.��.vڕ�r��?�^��`L�ر0Yat�������	�SXGI�v�rw�iM3ߡ�G�b @Oa�6�t3W���)[`~�o"7Yv`K^0(��5_�u�+�"O[0�-���O%B{BL3��"PX��g�ֹT��Q�_�ZȈ��� �̂���b���l�9>S�?BX������ؓӗv�?&�yh���]�Ϧp���>��=�e႔u(�iO����'H��@�d�~H~.�ܻ������'�����n��X��K��5�:SEs��:�3��m�IiCs�*�b�G�/p6�+��8S�?�^��X�Pe����?��	0��mg��N�n.-�YhU|�4|>̛*4=j���Æ�Dv��ޞ@Ӥ�|cHV��2�Z>���^_�x�:���
*S��p
ȈI��モ̎W�����r�03T�F�?Y�P��]��iq�|�J�M&ȉ�͋���r��_�pFm�+}f}�W�^e���St�?<|���lP���@�i�y�:��A�5%�Ƥ8�U�~�J��v
0���Ӗ�Cl�R$�XZ�\BH�y!�
��z�ڭ.�`g�r��p�Q|�2~�5`nFI����)�[y���p�.��U��ߤ�iF�� /�\-̘	���`�</bS�),������F\{�U��x�Wr$�����x�&���m�����:�����0��ԩE��c����jY@rjC,#��.u8ĪX�y�Jw��Y
��PƐk���kCx�Qڥ��D��hǗ��/�@�st����/'=�*�x�E�4ɉrvb�$�� �A+��QV�������?���;05�q��|D���`�ql�	Hm���]�z�B������U@I쟠���|N�$e|�Vcv#*��.s�y���������XX	 
��ף�V
���ŚD膑��⃕�C���=��tCmT�\�3������Q=`Ѐ���$ϣډ<�PI�Q�ə��r�[V4 �d���V���xQ�s9n��p��V?��-%wƻ
ܧ��gߢ�6�z:�j��OP���O�*���h�l�,��/��� ǿ_9�,���o�S"[������_h�;�k��E�t&FD~m�ԣ+���^"w$��!gB���/'���w!IB�C�)s_��2:�6\Ao�CUQ��|V��r�,���Q)
62�xn���E�Ռ����z�t�LR&#�P��ê��w2�~�q�z����i+�.ZqD��� (�FBd�(��@C��\��u��k?��w���띍�Uҭ0��cP���l��N�I|6UO�<�5�;'��J ������D�9t��9�s����>��8T����^$�U������0owc���ռ��g*0�ho����co�Qn#�(��[��)��59���]D"g�A6t#0h	�d�3=v����X^W�����>|�-��@�ɜ84c~S�'E���Ǚ�����R��Д썾����; �KWx����s��a�K�����l���}RgK�� z ��0])BN�����W����aV���5y��r��:ه��w��&�.�!e_,��tq�6�q[R8Lc�@�H���hD�sn��`*���4+�l=�b#v�h�ӊ��Ъ�2����[)I�����E������Yc+rt����}�覱*b׬�T�[8s�IK�ָ�e«�T���ϥz�'�c�J��$-)�Tq.�~R�L���ε��D�h��+�uCsL�'���^�8��Y�29�D{��+�o5Cp���%S���M>��m^|�QCQZ��v?nn���^�5���b��-��`�0��A3� �8v�0�?<�����G�{@ y�Q�cX&���pD�?ˋx�� "����z��8.t�4S���F�a�1�*����;�.9��(O�9���O��<���ѭb��l=m���>[��c*���B9�8&K
#O��G#�#��"�/� �h��E�^�X%������BX��#�	{N�˖�*��#^��-��E*k&*g����Os�a+�[�f�;+�2~�Ǉ!�¦�I��}� ȃTYlo�r�Ob7��]�v�m�5�˾�9�i�u�d�j]���������G�AEB������"����DO1��i�uߏAXa��]���u1�9i�b.����y�@��~`��5	��᥌p�[�2F^��p.�i�����ȁ��]��(ˁ"�Ά�|�99a�1��glf�Z����q]�*��s(�u�P5{�|R�D~�E\���{Dt�`T*m~ �,�U��u�J��b���f�w7�`��a�b�m�����>�K���Yj���1���6���]>�CngbT�$��_6"Lh�T�N��Q+X�란{B���\Z�9#���Ab��}&��aE��]PU4.TE���)P� -���ܶjHn����jy�h].�[G�j����7���[.�h�0|1~6��z�h	�$$:��7�[e�@�j�Ǖ(e��Y\�v��i7k��Z���PS�+��<h��N������D�g0L��I�X_���+�b�R��v����#�0�=�H���sO)�Qb���D��`�1Ff08��'qz	����Y-��#�AL����=5AuH3���]�l -O�U��Q����eŧ;MU�;��L�p�����WY�|�+S-��Lɩ����|SlI�"h�痭��ǜ����^+v����<w)Y9ܼuk�u^��cĳ�ٝK���T�lQ�c C�'C�U%zWcv��H
Ͼ���ꢔ�i<_��� EX����[/ƛu�������Hʮ��[K�K/V�	�-��ʩy����s@vK\��\��`�ZiOۓT��Bv�ӕ�T5KF��v�d좴�*b_G���E&|:
��+w��ElCqʘ�W?�#`��(Z�R�{q ����y˼���q�䎩�N������r���{a8A�m���L��9�,i��]�a0�z��dv_�vzv1L���hNt'E��)�JT�@qF�! :�@]���w��-�Z��፺:��%��	宻跳S�}�����K������Ϝ��ȡ�����x��8���=���r��n�,�Jt���*F�"�/H�bQy���s�ظuk[�W4R"�|�K��|�v���f��d������p����|��8�ܳ��1&�K��"�3�^'��_<��.������B���{Z[��ބ<:�,�e ��!��~H�h�T-A�@�Vw����Ryΰp���n��C�BTy�jԻĒ�CY��*�M��cLe�)*�1����(���Jy�����bI�LW}O�POw�d�o�����s��i��飛�΍���os��� .Q�_�_-���gO0D����!F��#�E�eG!����{tV^Ѿ��$�	sL�1)l$�vB}������:�k a
��X��ť��4��V��kK��/����?�3Ƒ,�;ݥ��d�R�MB�М%^%m��8V�V���Y�mwmW�pOs^<I����V�Tw��KA-�I�4;�z�����f弣Rn�u�Aw�qM^_Ǒ/B��h_�B�O�+ܜh����(���'�_�opd�'S��&��/  %tHD�jCpL�0Bj�Vv4���\�	Tt t�ov���O��R�R�U�ԛd���&0@+:�=b��bA�����ª =� �i��縋p�KV?xD:_���\2��QV:�x�Ng���DC��J��yEL�L��_�wƆ�������׸��C��K��rV��zNQ �>�P��i����JDN.��N��˯�p�PB�A�A�m��$k��	�}�����s�V�Iv��Ww��м��;�ɢ_�U�m��v��\`�vwQ*B�8E[Kz,��铼V�����t���~^"�bIT�Um��;j�q5Z{��6������M�4���`a0�p�(���� �0�!�x��v�2�{���L$Ax������7!J��Tأ)�}3l��a���i�{��k�s�Z��FQ^�<�q���h�9���jwOÔ�|^�[8Um� {g�G��@	�1�QY����e�ݜ��j.Mt���Ő�����'߳u�D��s���W<iI��;��CG��D�Z�_s��=�4c�� ����#��Cy0�k���=�Z�Ժ*E*�(h�ێ*������Mep梥�Ĩ���T�7?���GX�t��K�ecƆ�_���AEL��,��}��if�Z���T���m�lH�@w|�D;�Y}���}ۉ4Ty�C�N��+d��p�8A̗�t��y�
	�]���9z�h��]#:�|�j}����i�)��8>}6�7���E�Uƛ�R����PW:����2�#�'��F���Zô]���D��^�ϸ�U2�џ�!����¥�D�8�� ��c�xQ�{tE�wE�-����_�%��>X��c|�X��3�G��Z clT�	�H)�Yq¹z#�p��=B��{�G)PJ�)\�H�^ԃe����Sz��h�4�8.������{��&�0�h��<����E8�򏹛>?�0|��e���Ě@~o�Ps��(ľ:K���1_�_*���3���0 �Xw�H,��/���P�F|"�G�%'�W��Yp�&M��uq���C���a�GE�H�'����,V}.�Va�a����8Jl�ո`YY+���* ^ �8�a�"�2VN^ ����'�.�O"�K���r��E�d�[r"	����(���b�72�9��o(m������rԀk/n�J&:�xL�	�����	��_������ع����g�G���.�=ɀ���)+�E�z{��2��4���$��qޝ]���x�����(jR�nƘ�����j��6�e����VvG�������5)����ť5ѷ�yX���p�d��Gnws���	}���P�����P�H��r�������(���NC�?h�q��Ѵs�g��`��`�J1�)���Hof.��d�!�cG�?	�����@Gct�Y��\�Z'4���\͙��W�X�a��������g���#Ks���5���!�V���l3���r��s����W�`�gI+ׇ���.��s��6�%�i,L����Z�\n:�:��2��f�Q�/�m��k��Y���g�_�Q�m��Z��zKQ�|���ο	���qc�~���n�e���5~t���} ���%�e��V�9��y�[��4%���ZjEAe�5���(.j�O~ל�< ������%~�Ys�j �Q:㉬���Z �K)��ফxL��I�^w^i��u��J���͋`]0���>����%Uf���Lz!aSH���.DjP,��H�fփ"<O�sJ���9 �,}
�"��x6&_�Hi�`�K�;r���� Q8Ys��Λ�@��x2x�8�^�D��y/}�;kw�5%����
P��*�$Vn2��KY��]�-��)�W/$���;}���~�o\FY毮8��h���?�j�>o�Ut�,�n�)��L"�U����g?���R"����k���,&B�`�hm.A�,А��O�g������~�P��U"	d���GH� ��L�L �]�)�o�;*m�Ў&2g������Mǌ6ڢ�s��w�������*��~�J]/����KN�<f�V(lr�?4�e��`|���4~&�R�!�y(c�_0���8t<,_�,/���ڨߤ�wlu��8a�&�Ш��]q}�Z��C2��(A�`~PӒHX�֍Q�o��&�-�nU�n�T.H����I���yة�<ε��`��O�"i|�?'}�ɼs�*Z&���)ڊ�}���'bMu8Mt<[�� ��+��� m"϶0i��u���:Pϰ��'��)��m��wi�M���@jg��������F�	H�|R����c�S�=���p[84��S�ۊ�C�'����Ҧ2����W�.0+PQ����P�l���[�=#���푍��`ϣU[�n��N�)�~g�~	cy��z1�vi������R�n/y�[2<j��L�Δ����TC��t�� �n��i	�E��Mt��%��w����~e���A�CRU!����i`�\�5C&��Tk���R�VvP�u��G��v¶s�;�w�u�Ӌp�γ~EcXϭ6�5�p���A({T�+��K�p�3Nw�(�������=�+�Y.3*��殨�+�Q��@���WUi�F(�����JB��1Cgk��ur�G� Q#7h�E�|�!KRn_�M��]�$U�DJ��������v�S�=�y�xt�
�?��5z�ՠwL3�51��a� ���J���a�"#��-�u���ۡ��x�5��y[���u�|�y3�y��ukM*��8��8Gձ;��C!g
���)o��*0����1J���;��c1��/�����������WX�Ƹް�2?�{=�V{qy�$�F*kf�?���^�Uث��<�ZGI!)���~�'�����>M�����$:4]�-?Qm���W����'_��K��9Pm������(v��T^;n1#`i�>4��$��{���	�N�~�����'e�KI&��1>j*��A�����nˌ�S�0�%x��W�x���橣�5	����A�� ��'�B����R����8t�3X���1�Y�H�� �6�m��yE,����8��a���~��9���`�^nQڽ A���f��ni&�a�J����	I-��ۧ�Q�d��Su
������ &�t~w+�"�(�|�o�"��Wh`��1�D
��{�~|=�<�"�7�ϓ>�� ^���|��N���Ά�"�Us����������)��+*Nۂ�v�����`,do��p�{6�j�ꊲ�o"W�nt�6N�5qYU�u^{ɲi�[���ŵY/uw�=��T�eO:�X���L@� ���v�����6n�p�S9�ʪ�腩MkV������dfV��{�@��z��K�㡜4�fu3]b�G��X�'�EZȷ�i󮂤L���L���yg��R�3��~*�a#`t�_;o�E�=(�ӳ,㘬�B؇W��G��p1�_3%�c���J����+�ﳐ&oR֟r��bБ�_=�&@K���`r+cMZT�Sm1!�ؖ�P����7Li��/Iݻ�s/��͓�'ƅ�L'�7�P���U(K�����{�y�\�>�Y�P�wc��h�甴`Lf�k��w�q������p�j���5fNl#V%��,
B
�旯}�R�c�''��l�L�އ��y��Lh���L�ey�圴W�>A�t\�$�����֢Gi|:�|%��Ϧ�)�A����B�׍�Y���,1�nv��%3o�$P�=�Y���rv|ʱKF��}awl���Q{��G6�~pǽ���͏�3{����M�����&�J
�
�+:g".�@%��w��>;a>a0�p���p~����$X+�g��Y<�����0U[�aUC޾IS��WW�$h��NNz���H!̹,*�l�͊��hB����RBt¢>:Q�x=%힮�Yn�dmx��Kپ��ݧ	Nx���� �2�S[}|be�����8��d��_�� �@�j皳��	�I�kH荛q	kV��w	�QӫH�@�qpVWl����lgb�*�*�^W(ʖñ-��"F�wcxmC��s��7�o���F�����t�)�_^N�	�9���g�P1�J�%��%�/W�Ѕ�k�fݓ/��^�E�n���hϸ�/l&)�8�23������VV�!�;vm�·�����|�{��N�:C�����ݿ����k�{V�^�c4��1�A���t;O�Uڴw��o�hR.�">.�-a1�D�16��#��~�$�ڹM˂�*�y�f���[��*~]9c�����N�dƓJ+��:hT=4	�ח-�̏�)�adT&�"���Љ6��j�@�Gg��N㫯�Ӷ�+\�c�.Q����$�%�3r���V�_�}�{6�������D����͈�t�=��鼾#�|�q��|����8q��X�u�?0H��n.��{c�/j���+�j#��/��^���S��L�h4�6d>�-8��0��z�s�Z���.�޳����e3t�`}ǝ����@��rUa�1�-;7�
�(\Z�*�n�'�X�$��."rRL�AB Q��%1�|�#)��OZ��Hp�����!��ֽ�p��F8�Ơ4.������0p� ͇Xea��v��&�����o�x I�Y[��k|*����hΧoy��K���pů{���s�s9��%/U8E+BMp��g��!�2�|�'�J�\TR9w���v�S���@�_�+�ǄK����x󚺪\;�O�B� �X� �~ϕA�-���3���b�W{.$?n��~�\��)$���,��#o�h��t$+����﹚���f�n�� �H_� �ᓎ�L/2��8ٻ��>�h������\�<��7��	�	��q�� ��}�`�zl5�`�'�?;t|S�WE��i��A�Ȱ����@ӳVC�w|7�� ��{Y�زy�}�(Ԧۀ� 7�M�L����}�ܓCVl�{� k�)��q��ݓsY��P��eIR��LT�Ty��d����� O`Jd% :#�.���ԯ�6������5@i�H��C��,�}��TfҾ�
];X޾���G���_�(=U2��+�0M��a6��{*�Ȉb��L
����(�c��+Zi��]�_����"��^����۟{9o�l���1ު]8�$�8۸���l҃����~k�8�Q��iQ��Z��$�Om����(i(SudeK��(��N]̨уn���+s�K��h�"Mt���i���Z.�9s�Vĵ��\I�S�r#�ʉ�P ���^Od�/�t���\ؑ>��pn�;k�%3�kL},���<��u ��?|��sqr�9�u��eY�ޖ�X�����䃏�k\�"��{>Ã��k�G=�p�U����&zh"�O]M� �Џ�3�ⲣ����g�����0�� n*�
��t?_���Kjzn�T?6l��x��w�Y�A����:��MK	ØG��D~�i�˼�&|���i����2g�̼�2�J������� x���U0L,M=-8�=BN6�Zf�`b�J�C�h�}�2y]��?����ƣ�m��h&~��pmSm,iF.��:��t�U�����:i0֍J�;p���G��S��D���ʪg|�ƊK3R)2Q���s N�J�u��Nx�������;�VB@� �����Iep����)�J�eg�oO�Rغ+i��
�A}��KcD6JRR$8�#��mxQ Y\mv�E3��k^&���w<aYڠáT������D�����J�v(�\����eKY�&�y��w�|i7���]��Ũ9TDy���l.z�7UB,���F���K��#�J1{�"(��R��Ø�c]0�5�+��:����ԎUug��<ƴUZ_���@3�x�5,��&IGTX���VŤ$X|����zk� �k��4S��D��1�M�-�Z�|�Ե�*||��z|{uUmh�tRI��s��>pYo�-�7*���YP�m�m��9�0���D�;:��W�����W�s
�� E���Qiʸ���{�52D��5��p��~^��tn�⿽�*�VD/k��T�Ĥ(��A�Ir6&F��ǰ�(�y��,�G]�Bq��	�m��_C٬����!�'z��S�ϝ>f/�9���򡌸��dt�.(5�Ë#����t��>�G�(nS�4k� �ut|��n�rO�� ��[�񷻠����L(g��|��D	���&�zg)�Lf��v7r�(�8�Aѥ)������RZj)�)E�n
���Bϛj�Ž�{��ٿn����J� }Xw��`�D�ov{��
TZ(��'f�����]S�n�j+}-��oE}���6����7ޒzt�|u���!���o(|ȡ^�H���=(�gk����㰖Ɲ�L#�,_�_m�i���b9K.���x�"�E�����^)&܁�Aи�k���Ӵi��i�3bx��t)Q��j"�5ža����~�UU�.V�8	��$I�%!k�c�th�3����p��(�#����㣳���g/��C(��,OPܛ_���r��P��Z����v7�Ut��Ԭ2���WV�#=�۰:\?��30��:���gE�Xx���I` #�je8_��W����_Wn����[�������7�����+&)F���]2!���߬��E������(e=r�2���|eN��2q-@�`J�М~y��bB�d�EYA��t_e
xw/<\}*�4��-IN%J�Fz�l,�L'z�+�ղ��Y~�wb�ZJR�O�ǆ
 _��C�ut��]�"����"q�T	��U8#����Ѣ�hb+S�빻�?{��D�"��1G�9�V�Y�\�0���_���w>~�����y��EH捿վ��#��H�+��Dj�OE[p��3�*�7Q������5�E�	቙,,1��j�?�O��b�+|��6�2�t��]���������6�k���YK#�^��$
�)kh�z7�\6�����\v@���쌰4w��w�Om]|4<�4����`���R��3ma<{T#��a�nwB�n�Nm�B'fOr���<��nN{wPc8*d�4�@�����yMuF�lπ�x[����r�c	i��yw�xb`��Yw!�;�'���ŷb+�FG�c���g���Fw�k�Ŗ��L*�˭�W�<�������:�t�C�,qF:��4��)1㮄��Y���.�����X{!I�?��G*��UO�3Jd\p���KS��<�������"�x&�Fk-�G��_t
/�ʨa����c.�6n����/���6���a�0Q�z� ��T;v�J�};�Q ϩ�4�{_4��B1K$�7{�	�1>z�)�56�L�J�0��"�F��c����g�ӴR������V>?���e�xEy����yŎJ��D��'��t%�������9z�@��]^���� �2��Hp;w��KRT�Pc���{|�d��i�W��7q���9��Ɯ%��v���߀�4�a���H����î��7`��l*���)��	��!$�
�[�*����iP��>h�@�ׁ-}���_��}Cr���ݢW~I	�p��S�[�.�ʫ��.����1�M��r�)����F�v.�[6�u�f��!Ǳ��mK�b��c
@��/���2��Qs��C_���յv�>b�z`t̬������H���
2��J�&�Z�P�n�c��\இ;$�*��߯�?�C�*�+� �dۓ�t))˶{���J��Ze#��'�t�kN�*��� U��_���#�e��s`?�d��yi�T�ƍ]��g����P�X�V��V�C��������B�p!�m�0r��lI�Q�T4��1�!�K5�a%��q���c������l9�Yq<�R�J��X��E��O���T\���{�g)v*��gMԄ�42�����A�+ʅOhx�w�$;��6���g;Py�?�D�`S]F���_	N�p�D;9��F�!���1�Z�\�4�+����{����soKaTF��am�h���xɱ` "qy��ٱ���'��'ҽ��q��{G��v��E��VΗu���5�����w}��a,g����;�\*��o�/}�KHj��է���m$x����H"'T�,�U�@2��`ȃ��'��e)\����o���oP	�
��b���?x���Te�A�w��4�{��'9��<������剀2�]m�(I-�,�F@>���d��վ��x/�ߙd2������֥��#@��m��,ϔ����g�?N
�<���飏�'�
�����|V^��2�@�ȿ_�)t�t��b#?dj��	����g�Lf�����&fw�?�e�<<F^&=$�Ȟ��e�\�0b�d�,�^	U�$t3����ˠҹ9h9iq�Ie?��q���,�3=%��������zHw��������Q���>�9�wz��G��;�=��P���<�h�ٱ�N���J�uț&>��ɸE\u4�jV�آ��tzp �_3�vVI�����;���n(창:��.�\�c�뚐B	�<ۡZ%�a��S0�5�y�����S���O��$�6�^q�Zl)VR�OSU:F��t���V:�>���:a]��o��6��"Na��&���ę�E!�����,�tp)+6�b�Y�$ͼ�rŜ+L<�^+�pV����z؛�����"nYD�|����9}�JǗ��X�;x���R����Y��
�hJ���Q��ώ͋��Vq�Wc
%S�����ǣ����ǉ�k����bdR�MI�K�l���_�H��[�K�����l���y箮�J/mn���� �O�:�Z_C9�7G�0��J�(���P,i|�^��v%NZ>(��6>gsYP��,��s����YQE ��Y񻊱�mXc70;@�%����X꛴�@&��L4u*���������?���)׷bG������ڎ�'��,����o�f�w:���^�'`9^�˙�X�Lh# ���������T��1&S����VT��q�Y{������V8�$�@�f[��-�X��eF[�&�yln��bq�S��V@��Vk��`�K�8wzT��ҕ�~�E\M��0���� R*稚�ɂ
�bX�ۉ�_���d]�9�Ո�,`ȉ��A�����*���(�2��됃�o�)L����VW.�R_͔�lY`#}&@��
�R�����C����V5�xd9��d��FlP���~"1�#��0r�o(��Hj@�b
��#�e?cʲ�x���tp�?�c=�-�)�mcE�AI/08#JY����UBX*��f���v92Z]��鍫"܍|�M��p:`���M+�gj�����J�,$���PX��D���s���٫��n���>�C�@�G��f�|ZKrVD�m�����t��ym��(:h���#�;ċŌo7�G>��i.��t_��_��fPL���[�Ŋ�3��\?��N�����Z��r���UI�����x��D�g��s����5�Sl9XU��=89�D3�Ď���CX�\�*����i��<���#�J�)g� �[��q�mQb���|�={��=�|�(���n�Q����ך�<K�����؟�$��.L�U-�?ы^��D��˾y�D�s�j��+�����q�;�]�_q����P��hT�6��5R&X�R2�t@<3O��ܝ��8��e�b	���(����k��\V4��J�=p��Ej{B��1V ��pgl���ʕ$���Z�!��(_�'F���aXת3��d��u�����,��ah�����ۈ�$,g0�9kys���W �9ln�`$2����R�P�檄�É��"F��6����S��.�	:�މCP��:�''u�c�[�*�d�~4��d��GЧG��伤��\�`A�	�"0ِj��`�=`�o����N,�cV�M��Z+�`/�B�K`��y�M�G��f�^��N;,pָ ��f��|hH��D^z@u�X�����ƃ�ٖ��h̴<]d���m�^��nX���yYZ�Ӳ���>��U\�a���Tu-���WSP�+�N�L�1�sa�]5��Q��Ɵ�ن"��$����ܥ��R�+���Yǂ*�LA��]&�����0��U���w����eM���B�x����&�{;�%���؅� ��S�%=\�K�G$�X;��w��$�	8���k{gxĩh��i���wk����Go�z6���J�#�ȱ	�d�'܊�H�S���Cg�n/�g��O֠�ވ��R�%�K�+�8�/>f�hnrK�v���φn�C),.z��:'^�K0jۼ�'{ �m��3�^[Й�ͻ%eĂ�_��՚8�OEC��1D�x��k�7�4��,�v�L �ʿ�o�᤬�3J�z��'��2P���$��yW�~H�=�!�v���⓫�&3��!n�ȊJ@@�����=���/��8=�Md�?�-�7�cN7,>����cb��b}{��>_:�殘�L���qW��S���k��vrb�1��44��Y.S"E��o��+�u}���wˉ {Ùs"sǠ�o�t�������H q��q�vc�Q�QXH��D��f,j�{��[�}���+ ���WQ蟾|��F�v�,|��c��͛{�s� D~C0 �	XZ!���()r,�=��;�$<;.�.�|���٬�e)���.֞��Aļ�L�?�,��U���}�l��&��ؕvc-1�T^eu��ޗ,6��r��"�Pm{�h�@D>t��b32愣�y�`9�L`WCO�2RiU��%H�����4c��֡�PPpCCĲv]��@�]P��=���5Y�_'5zwC#H�;ʚNFN1.���Z^�R���5�^�mI�������J"�V�1�r��b���`w	!�l��y��x�v��ʒ9��/d���:�l�Q9�=Tm#����T�PU��X#�;�@�B���eO"�p	5� !	��HEd�EHx��T���!�[�A��o�V��=�\��U�� ����
(��Z$L#�#����v�� %FM�k�9��f�	b3�6�^��u�]�T�B�4�_W�����6hb�Ғ�'�Ha#�`P�)}	q�b�R`΁J�	��Ek]��	s�t4�kl0�R��΂�䛏�%��tV��WLV]!������?��ڷ�����I㦦���#M��m@�7�S�$[_�u��6�r'��J _�([���iA��0�IQ�B����8(5Yh��[�R���5��R���n�+�	��0�UGu������q��^��ظia�'���� :�%�+Lf�/��
3P�LО�����4m����4r<¡W�1�!d]�m��.;{d���X��p+E�c�Y�˸�H%g��h��=OpE�0b<zL���Hi��e+js3�ճ9DJ�'󍙸x5�����8�?���E����~G�r7
�^Aòr��v�>���k �=�h= _a���	t��{�߶a�'��Ԧ���u�B�{�9����I� )h�7+q7c��-�Į�)�t����sF�Kx��P.���]h��2��"c�Bb
2�/�R�t�7��O�����_%-"Z\�ȭki�2��o����K�FO a��2WW:�Z���>Nf�wr	0�O�s~�A�Ӟһ$�1y�/��e{��6�)���+'bތ����B*x���!�	���s��9��� Mw�J�cR��Vy��X�=L��)�VT1��7Jm�o�XCK���5��:�*'�*30�@���Q��w���|v�4U$��u.�[�+�y���?��a�@�>`�7���1�hy�3��*gx��A�g)��W�ʴ.�*5ʭ���ί��!g�3|�&��~
����W-���8	���'���L�Q�An�.W4���$E�'9V>���9D����BG�h�Dɒ���PPo��_t��g���<o�C��Yʾ��V�A�G{�ǵV�J:�r�S�f.��pJ1}o� �m��X��ۡXN�OK���nԫ�f��-�׷�V� k�v.g�l����hGP��Cks�s�SV�t��hwfe�K�T��yIeK�,_Ld�"�OC{往��PLa\��~�����r��A�/�b�dq�u�|�ʆ��
�N��2":7�ޜ�WJu��	w�Ÿ��������( _:�V�ۅN1���v�\�{��i�������8B鴞N��%^����*�Ѧ��XF8>X4�g��2O�!T
�B�
����)�K���wx3��x��ͧ�?6�ٕ�5� ��ڍ�t�.�a{�B*�J9<th��Cfѿ��,��n)�5p�lC~�˹/�>&�:�^�č�!�6>����4 W�A�!�RNP���R/+�f����=t�q���G]�\��	����ig58d�9@�$Η�!�f`Nx�7��JW[aY�SP�����F��Ղ��hV���� �fo �G�$���c���JBo�'����@��ۑ�*�ʨ��#_��fT�􀐟1>�<�y�}�h���؎�k�NB�\<��$;��[��GU��L���=���iP���dy� �.��*q0��Dج���� Wr�>�V��O���L����`��H^>�����O���ʬ� �0����z
��j�ݜ�ь�q+�����tA�W����zSչv�wd��`"gv�Kll�9�xq%>X��VX��ޖ�2�R��Q�S(yg��-��Dty�ދ���׿e��-���1�\xEl�$�4
�;�:`���P	ٜ&�Gg;��f@��A�]�x4m���a��#~�C�n��- 7�.�������h�����7)��U��?�I���z��r�˝�$6cͻʑ\{���V�h�����/{�So,J>�̧�M*�q�����	(��x��Z���]�B��iS�j�s�Υ���h6�AŚ�W�4k��.G�p���,�6����p;W |E��-�[�+��s�Z+R����oe�v��K?����G͊wu��Q#j��Q�KI�)CZ�:G�!IO����4�q�ow�s)��� �2�]�<c�R��j����4)
X�, ظh��I��z�.�br�דV���V#Y�Re'iU��;��G��}JHW�8C���z hj���&T�h�,��V���l����7��4����G	2��㭱Y�=�S5>�m ����5��3��♼P�g��:Ρ�A���2{:�}9�o�[c�eT޷�Y��B`ـ�PD��I�v;�.���� A�)���k�#�K�`Y{q0V1R�O~`��kG-����E�߿.:�g��@�uq��v�;�:Y�ٛp��P4"�0Ŋ7v��-�`b�AX�-��[��
-�*���'�g���}[�ڬq������鍰�A�h����B���k'����_ɪh#��L�NCX���@�М}ZW�(��v
�<uD�ڠ����z�w��vX�2	�%Yre�lF��v�K�w�5�J�gu���������=��!y��J�f���J�0i��[�@�MZ�h��"Y�ڇ��ν�=��D�����D���1H���]d�`HlWu5�{�c\Ҁԭ40V1�J����u�8n\4y�b}^f���z#�+�n
���^���<W������iFw a�h�d�!�T��Ы���/�nT@�3Jif��FYr����5;�*B^N)����8������ԙ�������f����
�1�����x!)IĲ�s���o|J�ZC,��ՙF�m���R�^h��~�w�L}�r#t'[�����_�Rk�b��uﶌ_WX�����S�3{Yɞ$}�mXߠ��J�3�	�s^��(��cyN��Ph�BRXHV�� �?}�u��o%�������ހ��K�:�p�7���tŨ\X�H_�B��|r�R�MvÇ�v�ZHO��[�:�$�g�'v�:^�Ut�����.��xOw�pOv׺��gH|^��ah�o�A��+�E�8B��[�~� ��hL��Gdˉ�P�ny�M�t=�d��F�d#�[���婘�u��jfd~Vp&����mƜߺDߟ}�|A׊�iA����i��xP`���6U��~�g[��]?�)�}�	�ജU)#�v32��~A��s���G"N�8��$���A�59�CIʣ�4e��@+�a�YOMD�����mؾ+q�N:Mf\�BCc�(�lB�6�A�n��XU�ۅ�8r�']hP,�aey�@o>]Fj1�;`����sX��I�l�)`�� =w���Kh%
&A?g���2R'���*<@y�p����7�1x�W�]_��[K����~`l`����[r�(�����"?�<W(�hY<(�O��0��)����&$zm�.��kF?���˧�I��� �j?��C½M�$�sU�l�����x��i�	j�w�HT��3W�yu`���|$���_}��l�S�!7�����`�Iu|س��	g"��]�Ur� �]��ż_����|$����#^$�^�F��թ����U
��ŏ�h޷�)�@9"Yߋ�&�G��K[�/�u�p��,�C�/��	�?47�?B�M2��t����>�b2�E�Υo��	�
���<k�n1a��{K�s�N
�va�B]u����ek�Uh՚�ơ�q�L��;*cQ����� +���+�~'N�h�&���X�U��7����h���/o��)3��M�� �v��˚�Ǳ �XC�'IgŌ1Sbt�#	q�8�~�6=@+k$2B�hI�9��`k���:u��t:�����:C��*�����K/0k��Đ(�W3qft��~���2��K6��N�j���~��#<�mk`�3"}�,�s 3���!=͌��`��\�;�\�V =F�Ԍ�t�(W!Fy��@��vZM�/T�{n���&���)OڕGL�|�?�l[eBc_�6^��<2h�&}�LD�ʃs����^5U�
ܡ��@o����Q�*�s0}�(�c�v�ӧOp�b{�v�c�	`����Ι�u��2����D��&�������TS=���kn�\�]dk�f����Iv7@�v���:���S|L�O����٣�s�Rc��\-�*�k������%SY��8���9���/�*��=�+��R����4T���5��Ֆ�r���k*����.�ݓrM�>&�[�E�������������;��8��|E�ۗ�x�!v�*�cJ��a���m9�ò-`~��a���A�H?7��y��� �y6ϳth�sTۄ+�آ��$Q��|�1���4 �?E�8��ys~.͚��� �߲Jjk��O�g}��)��#4/+�sP�o&<���(���]d�ԩO����^B� �.aFĵ���}��od#�F�K���u�|�����h��ld[�S�xf5��"�U�D��~H�WGD�G@df'�!����S �N7U����y��-�5��ˋ�Rk,{����`2Dڵ(��#hJ����@�<�=��L=��['��;̶0)����G؎��Z�KO�C�/��)KBmn��Îi�<����E�ب�� ihd*���'m�W�������"�Ś/��UM��������P;z QQl�s!����g"Ч�a����B`�)Cn�hfDo$xq�hD �7٥���b���Y��Ef��ZO���&9����>��st�lO���@������N��+D��M��P�F
�l������&���k���\�)Y{�[`5�X��I��占x���ٳ>��6S6$*��%�W)��- ]:t�#M���"L�ͬK\�;�%�Dx�;*��5�A֒��Vf �@(��_Y��Y�ۦ���95 ��,0FaՀ"�0�Mwr���3pu���-Yㆴ ����de�Ǹb4���ׄ�{�cN�遹Qerk���C�����g������?��5�. CL�<v̈P9O��ܴV��3�l`����_*������+�p����D��tR2�}��"����%:��5w�������\A�4cKg��}��}�|�=h�� ,>�X
2n�Q���	,�(�IRm#��oſ�:v���K6��a���j��iE*��|��ѐ�p�c�ݠT-��5��S�� ��h
D0f�S^�>��$� �%2f{^E��xE�(��ӒB$c;9�/����^��n���yݲ�J[��~��j6��/o�w�w�qCa)2��B�]˞���%Fd����e����s�`Ԅ�`nexx��H��ex=�k[�X���m_����M.�+C�x���[�p��!�M<b��*�m}�C�� �,G���nd�I��{�����X5����m���7ß\N�4��<_ܟ(;���,C�d7�ϒr�G�+� %R�A��q�%>�Ox���[��B�̚��# �cy�B:LQ�7�l�i�J�4K"v���j6���㓜�y$�-�^�׺C��L,�t��u��ݎUԉ��cz�����K�� <c�Ҍ	#�h�>.�����G`����x,�m��h�H����與�o����0����"��|�.0B�p����8�۔ڑ��';ܳ����n�&&�obӝX��ɣ��
�
�g����]J.0|'$�ۖ�q�[������T���6���ovH��Q�3ӌO+���v�/��'���y+��7~��&������VunVV��V^��w�GE����n���';x����1:�:p�L���G���IE�,	�1���ђ��܎&�2a3a_K�ȸQ�f�?�U��Q��b=�L����e���'��":�M�CF�Ȗ�K�5��D�\�'��2�zZK��e55���T�u���<m�ڭVgc1l[8���!/!��U��0����_EG��r�i��+f�y���t�O=�ʿs@3Bƌ�5�ƒ �Y��'��P`Վ��&���P�r��(mRt����R*�a�������b�~ �#S|L4�+�"�P�_/D"R����s�t��13���'\٫�`�AL�'���zB�U�7�J�Fj��	d������!Vد�9�'�pH(��������[dy��{]�Jj_!�Tma�W��g��b���mZ_BV`��1e�@r��]�l�z���n6�Eڲ.���ݑ$5�H=�F�f�z��E�?kW��$sJ���p=�E���̈́� ��Â��"v��q��E�F�o��{Ƙ�BdYctL��ғ��oF{�8XY��K!����	�GNn�;�<E�]�����)Ja�=�	]���1�|��]�uY.LU�wE��UV� TPQ�3amw�HUpp���-��/�k��М��}ej�ouD_5}}�\K���o��M��D��b���K������4Pi}G�~6E��kP��O'�7�_�v�3�`�����c�D�7Sfm{xE%ὢ/��G߯�E��k��ަJC����ѽw�uhʢƲ1�����2_��ڕuy��T�99�@����$�b���qJ�S�@5(չ=��a�j�܄+/��������H�>r6�E�N�eef���K��h�=����G���v���Kd����r����6?��s���Oŷ]���n$$��_�D�w�Y��s��q�7$P�d{��I��\������V �p���=�!E��6�Eƕo��A��1�~�)V�:7`!eH.eg�n�E.۱^q�DƆԦ�{�_r�+��8��|����h��2�$�'�?l6G���h�Nm���0����-���h6;�&zNkf\$�@~�놕ɟS�6�]���U�<��a,���~݄S��	�l0��]w2C���G�N�[xOWtsEy�Cm,���+�Ka��:���4�Zד�u�Ec��k��U�h>��0� S��lV���dC�rWs�vz H��es>�9��,,��XUh>RI�<O@$׏EH����7��
��
��"KK���aXծ����}���p:D�}���U�d��s��f�P���@��ius t���O���N7g���読�UP+���/&ԯS�ǋo�v��o4ʂ5ӧqGr�����ӭN+;:,��LHI��W�O�m=��uO��_}+�DNZ��4��oÙH�粿��q�A�!P&��mJE���)ճƕ��V+�[H�x�,�s06nǵ�Sf]���}nM^�M�hM̪���U��=�K�ɟ�LJ/H��d���s�7.��X�-��a��9Fk�c�Fiis�����<ʗ?ϏQ�&�pUS��`=��!�t�%��K�t�mi��}����X��ƄXp�˔I��ׁL!	֪�Z���
�Nyx���3l�:�ʭSPJ���R-�O|��靪��Vi��j�2r~Y�'v=:b
�$ ��{秭A�����4n�P̜<8��^t�� 4�@� +dA���с]L��l_$�<z�:w��D�k1�S�hrƯ�u��f�	uW�]�*�)7�[�ʭ�0��^W���@�����1̘�S��G�,�_�
�{�0E�gF��ml��d���,hd ��R/# ��pyO���=Fv�L\������#�W��vPPn��KP�R���77,���n7"#D(u�]��tՂ/�uFB��'�	�^#i�������*��x�I&�z$���K�m�	,d*,���?��!��0Tl0�ii���ƌ��K�=6�3P�6�� p�~�"�̩��v��������E��_�G��=݌��V
(��W�Yl��9�+.YW���8���D�%�nh� �ӓ�~�5��[^\c���)�:sį�m������9�'zp�xL��RNƪ0۷U�Mw�ɫ�/O� �92�g�hU�9O�JS��{�?�1�i�5�oF�f���4AfQ�׬ɧ�TXU P���Py��4
$�b�Y���/�����}(R�{=�u�>CT����������l)���	����]�Y$��+r�17b�h�$~�[N<>�ɧmRV��a�T�{htG�����9�a�N���슚p�ᵈ�kI�N5#I��e�o.J"�V2o�5�F?�}g��t"�_pU�-���RֺAWR68 �唪�#��۠���Y��2����Y�+ee�I��Z]Q�3_Ǐ�"��_V}�3!��tX:���8CP�=B6����K�	��sX�ya��	�V��u��U��R�M�W=y���bð?~����>_*���	&H��[�3�VX�!W���7�#�ƽ���֌P�l���1��/�ܹ�����W��d�c$qac�n
�~�+�t1�y�M�.���n@x��?����]}���^D�A#��&rlP��:��gʍЎ3��L�e�=����re�kaʽ�Oj����1P�+�I2tQ'�®wZJ8� �o�2k�A���n��]sX�P�}��⣇+Z&�]&�s�w�)[1<b1- �_9e�'��wV9�� \���v�m�Z�8q�3���þ��Ɲ{2j�"P@�z�~γˮ���v�d�m\��o�����i��1�k~��*�_�#"y"��v�\�JS�a�BR �~�҈R;?x�\88�V���N`��!�*>�Ǣ�����C߿�ю�g�fp0���e5̈�nL(�l�d�t�No�>u�ޘ�ZY[I����C�>�A�5`g�y|&]���{P� �O �+ ���>���9u�ձ?Ғ�*�$�<^�<���(40���uy�'��!�Î�;���+�,mGI.���|�oWŨ�Buɺ��O���u� �Y�0��ϴ_D��}��l3U��\d�,�jjrp�JV�'0�
�K_'��С^� ,Ls̪�C�yc>
�sD��s~����8N��������h�&L������JZ��՜�)�1�i$���㣗���T��K���a����0,e���OL^���c��/���P={O��L!�D�U[V��J{�������sF28�!
�؅k�͈��gP�
�M����P��|�(��qo��Jت3;w�-�O_S�=.'�~��b�hی�"�V����V
��� `i�c}rט�ȶ�P��	�VJ �;7��礏;.LA��5h�����K���|���<��f������w%�6ӵ_"�e���F�Ȭ	����S��I�=Q2!Q6���� ��̱XO�l
�F��
k4���z�݇�cL�`\�ꄝ5��h�.�,x{��J�w�K� _&��y�u�d����:���8�]wS�6�T:1������#DF�mf����6�XHH>t/3�2-CQ�+͉,L0:=�~���qB��mt��t6'�BEP�<��B�|V�v���pہ�J��"1��¿ȍ� ��N?�D~&�	ml1�`gcy��Ȏef ��t.�/#�;p�.rW�#E����� �Nbr\}��#[bgt^u"`���O}�KeA�:{X���4z��gO��`�29�~X��_ρF�pp����T'�İABsgit#%ߢ����u��f���;k.���4V`�����pK��t�X5�O�C�+�8��h	!���R�-r�#K$_L@c�Qu|�R�U�0�oN�ыs*e�ͰZ|��H�*��>!�ƈ&Қj 2L"�s;HqS���N;�1Y����Ǌ�`�Ca���\+�*�CN���r��]xwS���O�@@w��k"ݓ��	�^`5���y�-��jU��H������r�Iu7~�p�5�K��n�s/�k�vt�� �r�Z���:�Q,������=��#�Kذ�z�`��������h\WWFPo�/v�~���C!������1�/q�u��eH�__f3ae��{i�J��(3�7�ӺYei��[����G��I0�5;ɼ��M�ķ{�,h��*�X6�S/>��˛,[��y|Z_d�B�F�_�+��կ��Mef8�7�����(��/}���/%��_�$,�%�΃��uy�OTD_�dP���JV�v��q��2Kw���Ay�lg��	�j�{2J4y�MtN��˅��4\,6	~V�\՚�m��MX�"� a�\p�A94Q�s��ѩ�i �$����v��%��g�aP�H�B5�:��E*��ٚ��N>�#0�8}<��˘�B�,��-�$�7�T�"b�� ��?����>/N]8z��(!�!���f⒡��
�V��46�,e�eǁ�2yE������@O��/���r�����.O�z�"Т�]�����jm�v�G�qa'�iu�l%Y_6(��)<G����r i�V~�^A)���My�ź��b�0:��ȧ��lz�bѹ�	N9���XwK�O �ԁE
:T�ig�SLtW䶇�3|d�:ɶ��/X�>��YtJd�E��,B9"Z�>�\c�I` �� 8�)T���,��}�z�b���~�);�QT@B�Yk�/���#�Xt�[�F�f����^B� ƺ�O=���0f�:�	c�}�����k#��uJ�Ū��ҙK\�s�Q/����t�d$ª���R�[���p��l��u��}יsc?C���A:�	��ج|eKX���i��`�Y�	�s���].i�����(�`[�	'��׷f&��s�y���\�W���̄B���V�cEf��e�O ��F-��/EN#[2�1��� ��R���n���
zu�B��M���@��j���=p���A�t6B���;�)�}���1>�#V�>��:��S"m̉�	��{\�`iCӬN�P��%sǛ6a%ߋ�d!��5	�c�eQ��� �#��H�Vp�_�p��%����
�����{gT��P4;�<�Q����Hu\
̣�x)��h�7�y%���~Z¦-:�_ ��mBbMM��^#�d��,��C�-�*��	Ϙ�ۛc_ĚT͟��
���C��������DOgUDj$���me#I@1�ÁVQ��%�W�9�\ 	�PP ̻$1
��Mwh9�W�n�Μ�˚�T�.�qVO}��)����:ڱNڔm�A����H�6��^)Oc�P|��3G��7y���s@�0�[�1��$���,s�n�H;��������!`��=�P���H�$��ԡ��0�c�D�&W�b�f6>Ҕ�+��pߩ�q��ȼm���	�h������CH�:��e��ݩ���kn��z3}u!d�^?����HF��6�b�7?U���; 	u�>��)H������h��x�.� �p/-�	D}}�	E��v�G�q���̐�;��Z���ܠ���n�5��ȮX�owa��� �>i)j��3�퍽��<A#�)�,�]�q̋�Ev��"�t�Bڷ�8AT���a�MH�8�@y�F�?7יw+t�|@J���t������${�����6�#�}Z;W���b͎ Q��whO�`,}�����$�㮑 �M�.�%/�h��kfb�ΰ	$�L��r��7��P��J�CM�G\<O��o��~��T�T�Iε<W�<�Ȍ�s�÷s��������_�UJ[����s���/yq	Ng}��P�=\6�0d܊�:�a�y��K;��R�>��rgy$x	s�a�)�ig����:�9[��t5נ�d����.,�6���?�=��|��:ZeZ�/铺-��{Y�� ����]���u�C�f��`BO�eu���h8}��$�������G�<����}�e`㭼�W�7�5G�6��>�s�R^���z���~�sq�BR��<�q��@B�O5�V�b���}�UAU����j|���8�s��x� �y�����h�[�0&U��&�J����WA��VRF�3�kD�x3ј��nr}��א���]���\8��غ]T���ɲ~�`�A���y<�f�H@��Y*���Y���m���)Sp��%y�	Q)�wҏ�i�LF*s����
�
�)H��_	�USZ�0�qs�~w��F8a"sů���@¾�w:�
�&�XK:8$K��^w�)��ɳB�<�8zi4*������e7b�ײl�.��C4��6Nd%J�c
&�'xN�՜+G�gl��]%��"���(8n.�5����GQ�F��T6�j�>�ڐ��[&�Ύ�zγ��b��q^��J��z��)��#��m��X�-�Irg+�^�F��(u��X7��!��RTKB�~4��~�>^/o��ZpKU��2���}���۰!FY<�d�}Sj5��@��Y���΋��9x�g�4�ܵZHB[Ы��K�aƿX�C.�/mkG�`Ћ��迵s���<�=�����o}`�����;].:ѝ�}h4�_�q�p?�l�U�z���S�]�6KhM*[�L�txH8n~ȗ��K�r���3g��q:�Cbܘv���&�s��5.:���T+�y�)#��x�C"odT�F��ԡ�,�m���Z�5���[�TWb��h�#��E(:oAm`]��^Cm��/�!Zŋsac��x~��6]�|���z�4+�@��}%' `<�{��%UU�����i~>�f��Z�6X�D�� �JP;S�&<׍?}�l�P=0g�_F��
J� cJ��S�^
��nZ)ㅹpC�Bv@#����8OdrQ"��P(5�Ȫ�4B�q�p�n��ZV�:���.����+�T ��67�4V7bp�u�+��D�H&�:+i;u��pU G���8�i��֦�A�B=��ʞQo��'���J�D	�!��]��S�]1��(`�jޗV�#�M-�]㇒��;��ZRؑC�[e&r88O���"�x@�;��Ի��c����g�#'�����Ao�}j���ش��a�I�+�
1��|>粘�"/���3�����TMVQ�6�P��ͭ�Dڮ��mI�v� :����������s��*�4��S�H���>�y�D�)�<wF�v�3xO8��"��Z��☄� 
�9էew����H�����"�x���,��#L&�����H��A_���̠w�x $��� ���BX>~�d?��B�6�w��e�NdBSr"��5�q��r_�Av���	[��iD�FR�%7>/�-P�7+��˅��8n�F���������է��J�h(�CcM���pu��m�/TՏ{Z�-�.�t��vW�������1�5���#zN(�#`	�DCݍS�a&�T�����Q��C �c ����R���k�S��X��Q9�}�\��\�a��4ǲ�d3�F�/�e	ng����u�����i�V�.t�������,6k��aY�7ve�"k�T�� /�N���#�K�ԃ�����/N�?8'ұ�^sQ��MO��gȃ6+��76}״�%�8�J9��ܧo��ZYrN� �TH
���C.�c��j"`xa7�K�A�Q0B��
+ߑ;kC?�靪`��������St�����sAૢ��R��y�A˻]C�А�i~�(<�
�j�B�|B�0hm�)�w��3�
d�lq�}!s'��
��!i�~+��֎�� *�Ս 鳏�ݢ��"�<E������`c=��Z}M�B�~�Y���et\#"x�^�iovJ�� v��؀-uxOn��<��� %0�G��,E� Ҧ��1�R���ﯞ�yK�#�x<�ˮ:�4�^Xt��7O�>a��c��Z]b8�������D�lDD��+���&�^V��}�g}nL��!�F�l��1{Lg��u���|L�HFe���n>; l��խ��y�F�v�u�J ��k�P{���YI���#}֟߆��uG�K34��`3�����Z�d�����q�>�
�0�Z�%4��#��73�P��}�PtSv�1��m-�D+!�8�ش�XI��f�dfѤ�4/�٤�t�rq��	���V�]Z�[9<� �O #�x�����  �]���qǤě��f�/C�FBD�8-3����Y�\Өѩ���� ��M�����UV�w�.���{�����ބ"�i5��8����xȀ׉�a�!'WB���05E�J�g��^v3�w�=a��\H�U�Y���0IU&�(s�'.[Zp�:�tu�:ie�L{�]_Nc��!�u�%B��nހڟ#�0U!���c���b ^E�Ė��⫾'�uN�E�G�c_'���x�K�zr�rr�-�� �&�A'ٮ���[����� �:��1w���I0�|�O<�����������.k�Q���\K��'��g��G*7� ;�9��b7��,6f �(x���dZ&R~��[��6nTB������cl����v1��᱾��I��p�U:�~)�ؑ��_Bh%�-�Q���g�'���o�R���7���.n!=��Q;JlP�w0Y	�A^� Qa!3"��8-�c����H�v(�����78\c�jT�q��f\+(�#JvIH1���+Q����.S�4�� uL'}��Iyɢ_�u���Li����Q#y3�V�����8����w��t���yqr�o��&o�
<����w��<!?F�[�j���K'I��+YIn��6;F�V���>tp�
/�4=C )��d�SlJ�y ��7���(Ȭ3"21i���>ݓ]v�t��#��X����h��"hs�RC��(����;䲫W�:���� Uf��trJ�jl��ak��	�nـ���v�%5`m3-�`%�F�P�tz4���mt�R��uAOr�.	�Q�*:T�u[0K���̊��T�3&��*������-2m�Eep����
��ן[��e����ǌ��ETS�s"yb#_n���_%7;;0|��WHWcĚ���^�=�g��In�'�jp�9���F����Q:��S�)x��M��bn��a'#�XA�jz�L��)_����$:7R X�I�.��Uf��R3�c�t�Z�ow�h���_�u�/�*��@�(5�ǩ�$qP����]t&�K��q���@�� D��xǂ}g�#�fZJ���f�I?���k���-�S��t	�t�s��ڿ����� ;]!�eVk6W:I�B[�>�BX�h {����ME]�L�qe�	�G0�y��_�7���y^�"
)k�46��꡺��㭧��ᣒN���?F������H��qP5-�,l��($�v���9�խr�����0Am�\Cf�m�dqP:���% �HT�_)(���U纰Ƃ����kJ+#�C�7U��]2�����V]���<���'�U�q��V	A�FNY9�h	d�}�����-�MN�M�z�nE���e��З�')��Rv�J<Q�����I�TRd)�EgY���Ek�U��q��#{M�כq����Y��%��]��O�E�apج6�=*!E.|! =����4s��`����P�ҡvD1.�ʦ�PkxK�����霪��(����M�<�}p`����&W��A�(ǶXVmi&`�fP2����	o-��3�*8����%P�Yck��W�g/kD�m�*�)��z�O��wa'G������>�	?���,s&� 8���aFT��8Sk�W{0�c޺�������wX�����,k���xs�Rԇm�Ⱦ\�Ob�PKl�ȳ�������M���#6�	q��E;U�E����L�y�1���t;���?-h�����T��x&f��W�4ʿ�._r}2�d��)����L���8�%��'����E�s6�������bJR<1px��l;�gD�:��c�����ߕoZ���*k,�QדƦ�g�X�B�(�����ob�J����jϣ�Q����=�ma��c	�&��7�ß<;;װ�iA�/J�c :}����&/�l*�HK[�<8S����آ��?�D�ꝵҽS�r������:Մ^⯞���l�#j ��pI9 IQ�?g�t�r�]��p����"��� ����!��>��y��}}�biw`V���͊�n0ts���7�o�z2R$0(�aa���z��S �^˱vo�(�
�:k�6zY[ y�J���AH�j�QJ��*5����u�
��U��;A�O��@	�D���+���`�$���
�;�B���o8e+���D������	z�_CX�P�`�]م$4��neʔB��VN��h�eG���8�[e��u�KT�`���wL��>���Z2���Q�%Ĺ|e��S����v%6�R��]�=�3�Cv�9r��=�{�~:��;zV~P�F���=�!�A�[���a��$��Z�:���n�K�w�i���@p�����Ҽ��Wώ��q�Yާ!�)���f���+T<)>�1hMc�oK*�S<.����ɤyP![09�M�p��S�z���2z���6u[}h~��.�F(�57IxpM�4"y�9>oLYy�U�`-��F���Q��g;�uA�{v�TB#`UZ�T�tR�moN�`PjT}������R��裊�YF�ڡM�`�J��8 eO�-D�	/.W..�jUB�f����u�X��,bo�Ib�C��T@`������5J�����:T&�_��S��A⻜�C���"���8�5�,F����-@s�u��'3zi�KX��.��L��#8/�L/%y�(	�UiM.7}���[7F���w��ʇ��'3��q�!��3��}���� cW���VV���G���T�Av��2�����ᬙ��� Y�KD�M�Z���,3�����B�SE򽑽0�&�������W�n.Q�^��<)�!�X�%Mi2�q��%����@��O��vq���R��DIƴ+O𩇟�C�Ȁ�@����>��g,R�S�!����KU��PBA�����Z1�T�Q�WsT=��ex�@9Ź��z����g�FY��4hHQ4��|d���^�S�ϭ 9�P���k�Qi�~t�A����B�P@W��r������Ǖ�Ɵ}��>�C�,����C�lǡ�>P���w�I�f�R��@�X`'��u��a�N�,�. 4כĦon,W5�뫗�¡t�+�WGW-@��|����`1r�WԎ��[;�d�d�\��o��7�,c���wf����ߕ����Y��y̥�����Y���q��,z�XhD�~����77E�6��~c_g��ä8Ϲ��E�%7��3��o����ִn��l��b��se��F�1#?;�Z�����O6�/ސ_���%�T`�����eB�
�y�P38A`:D��{�G�i��u?췐ㄈ�޳�
ddHhu�T`�/C�K;�NbN�0V�������BER����^Sm�7��1:�Ak�7K�b�K���8o<͛�}�.���W!F��SR!,����u�H&Gq0�9�,�G������Ue]��m�ʫ;`������L�4�$�J�T[�ڛ#�)/?Jѫ;�m���������� )G�UZ<��V`�Qt2��h�KzT�4!��YN����;rK
	�KJ���#�-��A�AM�hOPUmO��@�Y�$N���]Z�ͻ��R$��=�7��&Ϟʪ���]�\�K%ܢN��	AA�5�뙢��F��^jD���@��*䏺�S�D�t�\�FO�:��t�'8a���f�8�*�a{H�ک�D��ũmjnk����M��-�H/p�71�2NT
���v!?�UȻ�8F;#�!�����NAMsdk8';ɨ�#y��[���wZ���tޣ$���@�`�[�2I�e8~��+�<��n?�<jkcԘ��Q*�OX�qc���
�@U�Z6R�φW?�iLkK�ر��n�s�H�{U?i��ږG�7�D�Į�?�q\u��f�tE�;[T4��6��;�"�e����1hY��ٗ��|���9~�զ%O@WA�>��#��s�"{mX��
�1ã뤌FM�����1خi�d�kp�s�.�+l���O�3�w�wR螠v|K��_�#@v��<~�ۄ�l��X�c����x(Q�.}�$�0,�ޤ�D����ao���H.M��5�(D�*qW��6��0���\�te*ma�2B���>g��EVn��ܵ�Y ����}��7��
J��G���ֳ��"���Z��*��4&�N��&Ra`y�h���C6t�hV��c{K�ҿ��j	qЋ*�h���k��5 �"����e�����< �o�����K4���X�V�
��Y4�5}p-�����*o�KV�T�(9�o���^����C�I- �x��n�mQ�!��O�b��+D����@91XÁ�!��i��7y�E R�$���ǣI�W����j�g�D�a�oR�|���å��jYMG�R`Z�ţ����,D�� ��I�$�[���㱣��O������B��G=����wFN��ɽ���E�8֢\p�"�H�ʾ�'�%�8hh���@�qI{���N�I� ���|m4c(����[pXnH0·`Pj7���QP�K��	��9�<��|�(������`�:�`a����T�����1��Y�c�I$���>�����O�Ć�3��P깶ʩ:���>����F�����W���&t�}W���䏨���L4��J���w	j+Xf/Z��C�$��uc����clJ��+P�����#W&�ھ[դ*V��W_C�/�dU�iT�"*a�iT�F��$���^�a���0�s��V��iG�1�@�< ���L�5�d�-TG,�0��j��_���O��BK]W�	¼�؉Q���S�s<��z����ĵ@��8\>���i<f��VFb�8�L���mKk~1�O�B�W��f#��#oG\��q..��G���J��5H��ۉPv�Z7:���=*Ê ֒Y�3S��"��OK?�Y��Ӧ���9S�η�8���8*6�����Xd@b��0'��fZOM��z�4>��߮���T��~J�x�z{��8񭷬jx4^@R��|yN��@�R��<��oD �u����C@�4��>�{ڠJ%ժ2.(�k=v������Ϟ�x㤃�ߓ��㉤,3i�9�ީ~��ٴ��2��$k�n�H��+7|������6#	[L&[�Vo�e9��mf�L����H(?����O�R>�V˶��0�'$�؉��o���M�3�Z;?�F�6�D<�nDN����.'Pi���O��H�c�i%�һ���f���[��|lU�<��_��!��p��5s����q�^��"4�����rY��{(y/��B�VA�2 2x��G�4m$IY���+�\ah���]�{���_�01��Q35l4Ա)��-:A�b�F59�?�$�oW�ĮʶFo,�^�`�#b�0�a�#& 4��Y�	��~硵�,d�X��h���H����&c\���e����M ܓ���!>e7�YHQ�A�=�~Ƿ�6��#O��I/�k|c2S�W�_�W�2_p�+T��k^�	R`�S&���Pd).�˅��Ye�z��n�9懺V����GApJ+�`,v=i5�LǼ?��HQ2���"膂��@^K�6.	�V��̑R8�����b6�'�c��+��\)�f��<�	�,�(���B��E<>T�Ae<��J-�����r��{ݓFMD6��l]n����Rk��7�c�˝��vx������;����^q|l��7��ݷ
]��j����i4�
}�����s�y��u�]볶�$w4�.!���yz�`D��B�*��?��@7���ZbUC��I���`����9W��'
*�����
Y�<���Ph3�ۻ��i#&13M���Zxr��f�+��#D2��7A^�8dOۧ��Y�zi��R6��ؠ��9�3P�%;4�
�O��֜�`K:|8<��~��q3�2�Ik\�M��Y�$�ZVI�F��	�H��w��")��q���
�䳻�K��j�і�s�U����7j2��\���[��h��I���=��wxVA6��?��K��g���[7��ɢ������(h�4y6�8��NLM,ᐮwf�����57Ծ��ZO����S:�C�:zT�������6�G���r���9�'�a���r�k��ʌ��#i�42�7B��Z�*�E���0T����*��e�gf�k�%G�=E˜������ײ�W	m�7���PY��/�!͠*��F����o���-��I�~��t{H����h�L>��"�Q��-��K|D���j�{_iա���IԎ�A䘴
�#F��P4�/_.!>���OF��$ :=�DK;�
�X�>z��Cآ�^"ݜ�7�Dj�����c'<��u:���j�k���D�O���\���u>"n���UtF�r�/���(�R���� ����]+�S+$U'���2u`C�|��m��5�:��K3���85b����W�{��%~z����?�h:���dr��a�.D#�����k;�oՉN��E�FG
�����]�v�^0`��?��K\O�]��U�}y�F���`��2��o���U��%�8Y�v�X/��j��a>s��8��xH5���"t��)
�����	�DU���A�A?i	VS��ԙ���t�����Բ���~����צ���}yN���zL�y��~q�&��)l�-/|o9 �!���I�(�W��������l�Z��b*�2dI���byt�Z6��>P��\��M�"�f�=o�iF���&GP��q�gs��N�,]�)���$�H�YX�"�|��Ni�k�,��^Ǘ�ęrQ�'b:�,�P�e�kZ�bb����N]�oPI)	�-^u��;O8�lm�ft(\����xྻvߙc���2v�n���'�D&�!�i�R~��p�a�g��E;a��O�7C���m\�+���.Y���B/��@�l�hM~S����W��x�_�C��S�Bʥ�C��4k��)�����[>�n�Bvᨈ#v2r�i��a���@�b�����k�|���RS�v��R��9��(& ���eJ�bn{�hۡ(X�5?Cg�b󧯥�;Ӂ.��%�h�����7�����M�Öf����	!���3AS��<#);~.�Ž Z4���#���#x�m�I����Wp�>_���8�\}5�HaU���.n��`���s��??=�_��E��O5@�e�>�r��}۱1Q��O���jlrz��6@�I�Q����l�s\�|_������]hu�
���Y�'9h�w'%mOc��="�s��R�v�S���!��~m/P�Z���T��l*1�����&��mt$�����AE��u�kz�(b����Pge�'�����)kwS-�c7��u��*�Ը{Qn�)t�^C���t0�h�Ti���0�Cu~l��B��R��3��m
�h�17b���:��kOc�����ZBg=�J�ei�_O�$��u�`x����'���=�����
tb$�@�a�x�4���ǵ�]fAf��:����[*�>6"���Tg(���B�� 7ᴉA��!�b7V���oA�g�}�s{��I�3����zH�Mx:#s�`J�Q P7���ǰ"�]�&�lw�{.�4	=%v^�:��w�(�5]2z���}c��M؅��NeF�	'$iL�3R�z�=�/GN>(������}�/����	��� �v��D%�e7��Zfb�oLR�z��+g��2��7��A�p�;n�OM�O����}8�A����T�C��e�	����dx�-yZ��n�:�a(~U	�!�N�ۮf�o�S��/��o����W�"+*�D��U��G��6���J�1�c_f�y�^����PY�*�In>S <�.Dg�7��V�Q%|~���Я�]�
t�^3�\��h��6����Cz(s^e[q(��&
)�~@RȌ+�w�#ڄ��g���ߗHERh�{�1&���� {dί���&Khw�moj�nuE��\]����AK���cX~���xZ�5r�y���-�]�=>?Of/vѸ���>�	�@�h�/�M�k��GӃ|�	�Q�(xЭ�߻��Q���#��G�5���sC�%1�4_j�?�ؒ�h0B@�?C�
�z0�����Z���k�1o��$R����a{�o�}V!x\�@ǿ_�&�xʧ!G��o���U�CV���_�ë��߇7���"�A�=�����o��_�tli.=�d�3���7'�0(N��~�\�ƽ�j�u�~zhTK0�9(�U���=M��"�s�Ss-b�/ɦ�i��5����T�zt��kS)�9�]�h&h��(����apO�pQЇW���&D��Y���=Q�%;(�fw���6��Ŧ�+M�T�.3D5��Ρ�U ����D�ox'U6sj�&䅣<`��,
�s p�d�PE~L">�d�yxI�|3٣�7�KK�La*� �묦�<\�KM�6�j�˙~�*q,�>:���[�� �IB��$��Z�4+ϵ�����d�n-�E	اn��WJde(z�a^�;	\3~щ����W L�wfY�J	��a���y��>���p,���7��-�	��V�	  %�"��"����%`�q�쇆�n��YՄ;�{��3���V�m�����fM��t��Z�ͳG�$ 2z'��e��
�qA���\��KDt&M\+8�&�d���ĔIg�3�J�DwDP
����c�g[vs�۔:����h�,�kT�]�9e/;+��W5�&Qmok����@����C����B��0��1��՚�l�n
��N��9�#LE��D��vJCu��ҝ@���.�P�:e?;TA�`v��a��:��!�O�:+��\��D5�3�qo�"��1 H9p?Oht�X�ϝ�&��/�n�)6���CY�����E�K�^h?��H.�7����WT�0����6x*@h�Z6|u���9c�/ℯ��EK�QY�ޣ�]���@���a�LG���W˕�F��Xz�{S�(��J���(`E�p��:��z��Al�EKHn���D�hD���������T2�瞣��]{�����Ǭ����g�2�A���I}�p�M2�XD	f�6;ł]f]JT+˧w��'0�A�$��a��W*��q<.R�Z����Q!	C|��@����l���}+�$y�����B��|-�2;�X���;W���th#��[�t<�} X��·K���w��IU�:��O���u_�	��J�:-f�(�I3m�	��t|x��ļ�F�o��!�]�&�6�"J�sT~�����y��C2���R��ue�f��
~�دDʡ�\��zS���
���x�>8����a�Þ�����[輆���ib.��a�v�FU]��`72]�I5�2�(ձO�8���rW��BkM���f��B�?�.>��*�H2��� ������f��� ���F��B'�h?��]m�(���?������ا_\v�v���*���S���b-Qٗ���z��0l S0[*��%lʑ��V��'Qfg�눵CY`Ԍ�c�E�B6:��#�=ʫ'�H�]۲d��P5p�b��9�y?_�U|I�.���Sq� 8!ɋ���^V����Y�c�n����'`wҳ�U���An1�Ee�v��8 ]�+���~#����Q�?mWXւ��`�����P|�ߓ,1��ܿ��Ѽ7��s_WR�Gș̻5E�țpf�˛f�з��ռa��0ܑ�ٶLؓ˵[��(���:$2����/�I?�S�
j�)&�wc쀬)�w��K���u&�RAitsP�˃�ǎ���>��O���K�=���B��I��ּ�<CU��o�1��1�T����u��� ޫ�?�BegM ���e�L�m'�n@/�CϙR�VUH��Ը��\4y	��+��A�m��l8I2�����M0λ����x�u��?�����}�J��/�..����"�.���wqjq�xFc�����* �X�;�E���9�����Zn�)xUfp�n�զ7����U��x;u)	��ā�բ��������Q���_�]�=� �P��׸Bg�J��5�)��F���8Қ�6���'�V�4�?���t��x��ٌ�v��[�� �����uPD9i-e/� �}ɂ��_�(����^������v|�����#�_�c�s��t�7'���U3�������{}������i��;�r���.�� ���(���E�m�t�w��|�N�a+�:��'�A��|S��+�/Z��P�V�0�	W���{�Q�:д��?/��r_��M���0D18b◇D��"젭�75�K�e%��S-i�����Z؆qn�h��%`�~����T�Y�s���VR���QR!��R	M�6�"�qG�²� ��K�[��4�W�]vD@d��[a�m�]�f߱C����,>2ѳoA̮��X�,O�!u�f�IB�E�����g
��<
��"箳�����y��7�@@`�����*++�b���7|+�U�)W�4G?2~����J4/�]�����y\��+�m䕅�f�,�1Um�tbM2�E�Z���`%Ef�V�K<�����a�G�.�r�A�Þ'����"�D�ѥ�yC�m&��r��؞��`1}6��m��צCvz���O�=�[�>oJ�O�ӧQ�zQ��������G��M8����k��`��E� ��oAK�<�e>�����*(���4UJ刁��wd#�M(�߾�?=̲�U��8����	?IA�V����4Ǔ��v����;�Q͔;^~�p��i�7�}���zI��}j��^R3m�@F�2TJE���x!�w���g�mמdѓ��?t"�R+v=؏����cgˢb���gbSf�%`!�OͶ_ݴ(�!Ϝ׾�
��S:]�M�	��+��mb�����R5ٹX���fdJ�j�F=If�G�*�g�%bmD"ۭ���mN�N��f��&tǬ��,h�N]<3�͍�@�vH�I��x���3KKyCDJO���;��z�jUQypZ�KM$�G�M�Tc��:����Df"��a��Y
Sɓ@�}Jc9aBj��ȣ$�{&7���/�r���Z=�6bhs 8��8�mۆ�3^Dкq� F_[�*�j;BQj�-�=��D�|!:�Qv��OK1Ai1�-^a�ޖN�޹G]�/g,%6Z�\�y;g�8���^��-ޙX�z_t��6�R�?��ꀯ��%��V2�x1MkT�4�C�3xP?\	Z=Sv!��<9�T*�0�����Q�����E_Jt�����ч5�A�g�@J��(��w̠(�0d�=�)��]�m����~5��tX��/ۅ�˻�h 	"L���~!s��!^�-�yI^�z�����X����Y+�H��B�r���;uӥU3e�)cm+�K�1�0�񦕸��_*��3�#�!߫��4ItpA�!�y��5�f�=Gȑ�py�V�\��$IK�#��vtL�8�E �YBq�؄�<!*{�v�������?�������ǅ�G�n�ݐ��s5kV�s��f�����o�������I�9�K-}��k�?������7���.HN�%��c�a��vL��$�
�=�?��wRp]]����놐v ��Ua�H���r���;视;��
��~�08��e�z����S;�L��p4q���P��
�1ܨ��>���#��X���p��Մ�8�a>��Q������L6�1_�Xqw���0�)��X�~e]8��.[�Rʣ�Z�p�!�O���X���~�rY,RV�of���H�Ìu~��5��t3~�?���_�=���\�/7}a�W��A�~�R����"J�!-�� �D��:I:��ޡ$p��֜��j�/��0K��б�@�IXE�Q����pY�^w��"M�7�������e]���%�!������P�z�֪X1{�4�M����[,k��Y��4d	4l�L]��$I�Qӿ��N��7D�Z�v���uy�R0�<VSev�Tf�}��Bb`�g�!4��̲�*vHYco@�d�V����7T5�5�9I�3���WC90p}^苮C;�Xm�f�.H��AJ�|Vb�zxS���"`3�M%�5~�&D��"ш�XU�Ϫ4�'A�!VL��X_�6	'���N+4�w�j��dvXHz�N�k:{$�Q�������.�p++͑^L0b-��D�e:�h��Bá�t1F&�A���ċ�x��p#N��(�@:2�9���s4&���נCޡnf���"ݍ�JZ�~v�8�e�_��� ݈8��=W�d��;�PKV���	q���	?�=����snA ��<cye��ɟ�G�cp�3(Y�0*�D�Xl�oٹ�_���+�^�U���uq����}��5£��W(�^,����*��N�\nJ����Z�(ߦC��_�QPh��Ȥ�DP"�l�ѥ���Ic�=�{npA��-�$�R{�����,��2\>{͟� ]�I��3Y�ٓ�D���"9ta����-����؆ΉWw��T/G�JYg
w��X�&'$�\���ݱ��@��Є���^_K�5��E�+��9��Z�bZ���:C���Ӭua�W~P-�^Hr���c��/�C�/?�J86�$�� c����@ݰ�����H�2����ʥ�C�D	�x�A�^$Y�J�P�<N	�@
e�b�9Z�TD� Ƃ��!�Is>�c<��􄒾���|sW��k
�5��.ǃ�mh��Կ�.���V4�"���9	PJ��|����W
[��k���F�#�>�8?���!4�����Q `x�ω:-���:�ר h����>�L�:��ق�� ��&<����.�URcV�nh�`p-O���e�є�`P�)���@�y.D?��مmD�M��}Y�ơ^�%�!��,VJJs�@����ŨN��ס�|�n˗�;���˦�jjE����ϟ���Q2���ոp3Կ�Z;�Y���$����˧���;��I�� z�>ᨴ�����i�����I��Q�A�3�v���rG�����d��Q����UFf�g=JAu��`-�t"h��Q$��9B�p�6)�뙉r�9�������|���һp�<��7��Ԇ�؁��!-��ȂUb�\�h�@�66�y���n�7!}��^���L=�ǝ]��+h��ķyb		��ڏ�R��9?l>r�PVZ2�������t��Gc�¯d�J(�Ŝ�BP�]�z��V����չ�����r/#�o^�~'c�����M,���(Һr��|͹�I�в�Z9��.�t�9_��&�q���pS	�M}J*9|t�C�tx˙���[�.:��;d�_�&�=��5�+�����A�Elo������k;���B@�N���/��Ў%�͒���m�l��"�b��'�8r��;K^����?{�x���Kd�ĭ8Y^N"#�Gp�H�'᭭�,"  ��y��KNzrO=N�fD��k��bC��*Y�IIp�bk͔�nd�K�xG^���EW�60 "%$F��T�jF�c�5����i|�%GM��<���C������'b���/��NCY��j�<���k>uLK��&x�=9�Y���T^ҩ��S=�=N���p���4ZѸ}`a:-�W�4�ae/e�J��F�i�xϖ��CR��BM��d��KńUS��!�A)���ߥ;϶1,�p���q��݊["35�F&|�)&7��)\I7�a��xı�e�>w|���Za����A����"{��|G�A�=�3'�*/�1��#�H��'��xP�g��*��bCRUB��K&z=���l�@Jd�u 7Qb�9��N�.]-��wM4�����^�Y�WPx�s��<C���%(c�y�U�BȷO��p��e�p�T�W;��D?�ӗ5(tpE�=���Ʋ����wѬ�y69� ��*R�ƛ�l5r��)�S�W��5��0w��q̲#	��Mb���Ü�׮���+�w���KʕW�����ߵ??(�h�����c�#OWh��|VN(x�e�`����=�b��ad���3H��G�� �2����cdP?{��s�m6m	�}����7�6\��~��G	����gG}��8(���p-�ܒͦ�ƽ��ĸwki/~�F���Y(?Y�ZN�*�?��K��M �H���?6t	)ў�����5hm*�¡U��hF`?V����;���Qe��,)[\��-�F7;�3�l.�{��e�6�����L�?����]��Ƌ�ޕ�),t��i؍��U@[S�2���9���l.фx~$?B��C'a�oQ
�}>;���\Ȍ��5%�pm�{f�pg���ͽ�_50q ;Q��p���.ٛ�zg�H@�t׋}��Q ;p�Ri���-I����(c
.I}���~��j!� ��1C��P���9|�
�Q���_��nYa{�{GH��(1~R�X�)?v_b�lyS7<��|�-1�=맜�$��HS G�ǲ�2#H��~vb��Lz�tp*�
�Id�K��b<�Y�v�g��?.8����G�}�u1��F(�3�3�Fr~O��6�.)e���7���͊Hȇ�����Gc;�Yf7�(	V؈d�aw����,B�h�$M��Î�.a���LQe�|L0��z;�1<M����J�-�`��j���e˾�C�~dJ�G�O�k◥`�pHd =�l[��� k���l8���M�������D��'�X7��=v`����[P��Jd�[��I�A�h�q�u�k�gu�N���i��Wk�\�d����{#�o��V����o��*�&dst�E��I���9?�ԸZ&@/Oit�R�����2+	^-p�/xL�ƿ��"�T�rA�t�����+E��k�k�EM�3�M�W��+��DD	��+J	�ע���0%dɹ�ޯ�E�tb%c������~>z�t�ײ�S��Ձd'omR�H� ������}/�pt�`�o�����*�L��$Dѥ�B�Y;f{zo^�䐨|���C3D����6=5k��!��8��V���pt�5Zq�rם!r��ͮ ��0������Ґ{~P�@{��gXSq�=����6Ej�������H��ǐ�o�(���N�X%���
_9����Y�I���+�ё^_T6C�%\|`��ڣ^�ϩٙ"�ݏK]�?J���U�<E��՛��E�����#T�a�Y�h�IYkBt ��;��6������N�/1<)�����+ ��rM/wF涊{�'riҕ���
ȵ�J�js�)Ե�^��[>�����o����@��x,��g�M�6X�6��ߋZwW�!i����jt�x�N�}�._���ِӆ���H��t͜
n/x����tQv��*����R���^F���5�ycK>�;��'���s�E�ԍf�ϜM���f�&o��h8 \&��]C�S�A����jƆ����uB��	��|���K��zi�:l�o�(Y�)�F��@�<q
1�ka�n�*~����
rq�}.x�����v�@1����:W�5�����V1�v��ϲ���xvb���?"̀Ī1�,ڣ& ��iZ��Q�q�B]݇��.`��?.�h�Tf�7�M�f�C���'!��jL�L:��c �.�]r����p�۵�"1����촫��0��t:>��{]i$�h�3)v뵿|�q!�O5��:>"��~�<������4T��?����ަd<Z�d����L��ofZN݊�܈ς�����."�K�O?F�v�Yy҃sUNl���ș�y��ݗ�dvY�5�!C�.�dv��D~)�O�(�,�!�U�Ö��!ϼ����>���徏ԥ�<a|^��'v��� �{�c�6�������q�d���7��!r��fzQcP�R�f�$N���O\�gdQ�gL!�~<�#�������#H!P���K��Fëֈ/V��ډ�z���aa,˚�ڥ$qE��н[ݺ�PU�.M s7�t=�<%h����A�caدgiM��]�������2"� II�{�j�L�%�u3+q�:MO1�rM�5��K�[�	L����_�Гe�RIcbԗ (%V�q��_���n'h���'���ַ�[0R}��T#���ѥ��θ����|'����݅F.o�Z�Ǐ��Ki��@FE\���s��'LhF�=C?�U�a����ݤ�!t�Sq���Έ�[4�X�,;7F!����1�g���|ױ�˕�?ߍt�&�Zs�	�
%L�5���N|�iP����Ɣl���Y��|�	"�MSi�[�v�z�H�#���W1u��n{�M95B�^&%t�f⶝l֧%"`�M�z����TQDy������A� 5�DAƣ�8��/B7KC?����CC�����W|��=�e���Tb��*)H���6T��NNk[};	��{�D��ܧ7�������mŽ�fB�(;�C�u)氠mo�d+�y�=���%2�O��=k�$�5Z�Tk�Fm��PH��k�uRUŬ��T�л$�/�D��R����#�`�S��� h�ɬI�̓�;�l��9�e ��+xdptr�	E���ұ��'��|q[#��'%���L�����=ۜ����Gg��������O��Iv�4���` -��,��0�T1�ۯ�ך�W}v��`C||�DH�2�`��b���:�������m�7��5w ���f�1Ir��\'&1b�a�1��|xDY#<���B�y�_�ѽ�-��O�R��(c��s�Ġ�H�-�k��Q7	L���'��ͽ��E���{H7�Ô/�E`��J��f�QE�Huy*����?�6T"C_��'�o�j�K/i����+p��27^���r�p���s�*���ѽ�톾��@А�”���-�'~�M������Jjx�A�̊��_Db����F���fP��nG*B��Wu��u�D ����}Þ��;���<� �B���	���.������!�����άIpn��z-�&LK&9/+��uYb٭x`[x[��e�j~�<\���A��zT�i1�t`V͌���Eek�{ǳ��س�����>T��+��
O�w�J��>��hX��n\�H��U�R�ۅ=Wk��UG�:��Et9��)2ex ��˪go.$)l���#�n0��������`	�[*���fb�,�Y��)�����].�*�xg����)���e&�2������2]%_dF� ���'a���0��������KLl�ꗵ�I�W��eE��ddw��J����;��>@9R�$*��S�'ri���Ɂ㸩����aU�y ��̋!�*J�6���(>�y���67y6�EeJ<j��&Ka5/���!V��lf
F��lFE���~�p��-f�a����n�=l-⁊C8`��Gz�#��������7��0����f�>o�U�������zu�D��6P�x���f�'*ʗ�V���R�|R�	����%���Tw���v���xr�h9l�{��� ��ӟ�O���RZ���J�"	>�+A��6���U�!�n�Y����ɏ^�)!v�"���X�f5"�<���-�/utB��<`}G�WK����pV�6�9�#�EY��1��D���2s���5l��sz�ľ���ҷ��r�RՅ#�^6�B�8S~T7"E�,oC#]Ծ��1������!�SE�:���4���.A{�X��5}Y�_5C��#?S�]��:y���1 9�B�"�ޢ��;t�+?�z��;�f�[t8�mȗ-�6W��h�_B(���1uY�t�T3�����4^�]"]�����L���X�]%Uq�.qg�m^����6ݳe�9��\%���X��y�����2��C�v���3�zz���z������C~Z6-���%�'E�UIaU%�x��t��8wL*��(V����g�0V����y�,M[O
oMn[��.H(�`t����}�-��w�g�J=��ff������S�iLU%��	gk�4���1ƱR�Q3}��E�i�n1R��Dy�@��'�����RGd7zMx��tF q�#���`ٙ���gE����ޞ؜�z1=N�p&��Cc���ޣ�aGx��S�xN��a<���Ժ��TAY�S ����9�@=�LU1��Z�B[�ݲ=�ȲE��S�r)s6�-Q�+N��zD�vHө	.\/�|Ʈ�"�дԑ$Q���B��2�k�o��V���N+��U̞D���@cy�=5���]��n�m���r;	e�M���)è�5{�0��L��U&狼�G�v��-H�����yC�`~I��a�<��}ޒ��F�Ñ���l*�s���*aWB����;FT7��2R_lƗix;�\W�:���k�9�F2A� �OP��t����[�*�(\�O��x_��E��*������I�����Fj�e�a�9�� �P����,2<����b=� ���lP�)����fL<�A9��?s`��o����$a���.�_byO��q��Vԏ�����_\��������6n-�j+�Y��� h�zޙ� ?tA��*@��������[�
-���0������w�w�ӛ�����Y�����TyE,�Ѭ3�X�B�`u�$�@宣v���\k��ڼ�F����r��(���>as䛆`�b�?&ʆ�	�UQ�t�ޤ�@�%.�1�7�ҿ����$
L���Y/V�n..�a����
�s�1��)���
�'��"�	��c��G��څ�+`����|��<7�)�E������s�Û��m�i��H p=��xq:����[�!��~����2��?1�ż�e�K�Y�- Y�9��<E���T�%O˟iIʱs]h�T!r"�	����*�ӝ3����ç���5�ci�9�)�%]�3�]�z����DԮ��L(T�%p�z�G�����<<�hB4Q�����i����n�Ro�(�Mw���CK|V8��^Q6�W1C��,hNy��ኩ��n���X׾{�$K�-+XR���
zD�&8���]��@��4c�n�Y���1��ŠF7�8w��w,�����r�����\�� �R���o40�rL��v5��ᠾjU{��{m��=���u�b�=�Q�����R�5䗲�%'��>��f@�mO�*[� ȵO��Q,B��ab2���,�^Jt�,w�
�h�\^x�s��AT�AZ�A�e����DB�,��qH�?í۶�ƨ�v���Bk��ub�����sG���Yy{ v�Q�9oA�g.�0BTC}�Hh�UX�g�Ad��n�mA�Q�K4a��>��^k4��o?y!~#�	W.	�(� ���L8eB��|s�����1c�1�51�%��B�YJ��ǈy�o�B�2��͏��������[&*��q����b><�#�ϻ��d��Y��v� .�)�-��E�}�0s�H�S}P�`~�N��FAl?	��o�V$��"�3k|;�� n�D�)%���g��
=K!�_��Nx��&Й��Y`����'O�󔆜 �i��stf��Ɵ&�Q��z�qq@��^t�5^k�~O\ҏy�����H������y8�HGs)�E�FC���V��99�I@�~s l����s�'<�>��g�%XĶԟxJ�l�#�*6�O��`	�<�m�M�Cءʅ�;�Y��i�v�CB4�\7��*� �S�W
�.ۮ$l�MŦ�y�.�V�H]��z�@v��G'aý,���}B����s��E��>>��e�n�w�[:���s�������+<`��Y(A��O�
B�)at|*h^xUOLk���#�ܸ���8$���(�ig������l?>|W�37+�y2�!��{F�t,H��.��_�]e�T�+D�28��5�]xF�gq!�RL�5�\&�K�p�'��Vϗ�"�|��3��aP���(��vͥԲ��LCzX��Ey������
Ñ�89�  yCI?X�����,Gts9����Z����)_��j�ڽٿW��h�*k�-����	� �Վ�x�l��#�4}����J!Nᶦ��y�
\q2b0�z�m̀�pyo{yD�,���x�R��e��Z�GE��\H��]��mC��ቻ&��b�2um�� ݤ;�� ���  ���bJA��t�$�cA��C���~�E �'����
{>��!����O^N���a*������P �.v ��_� n�����r��
�s�Ş脂�}�n�f�\/$]���1 {��K��s�x��AO�V�����/�N	����MO�+c.�}.��I��{�|��n=ąW��
�;!��A�����
�ws`�jW�n�K�^ by�y����dn�����W��1Y<�,�޳��q۱��G�0�=g�߅�i!K���/�� V�O����Ὸ`����t�|)y7���{�Hڧ�3IŘx�N����5�?л��5��O��y\I�n��v��b&���6��Q��7���=햶<j�.zS*�jh�cС�RJ5��yr��hZ�.��@������+�2ށ���)CX��'鸟I�wI��n1����g�͖~8���)��*s�m��q9xO�彞��:�1�]����{9�*����.��7MQ����iT�5��Ww6O���a�<)��f%X,a/ʙ�]��&��3�n3e/���kk��
IhF�����U��ô�JyE���;�=z���� a>��	��8�ngD '�&C�(G��-��I@��>�=z^_6� ���2�������L(�P��vN��_�(Z�&$��������2�$�K�4N	�N�z�R5�`m�aŎ���س6�ЍU�Xsf]�F��N���k��E�������r{�儈����s(�|mbVRs�#�w`d�GW�}d�ͱ�#V��6�y�����ӕ����i2�`=��������zaؼp0�)�6	Z��^I������9g��g�>�r3�l�����[l����[��� m���Ko��3���9K��zE�/��=ji\�$H��D���^ ���7&�Fc�^�%Yg�G��k��|v����OvI��hd��ǳ`�*�<87��.:� �u����>83��}k�4�s	C ����X3v]�����@�����!>��HB����Z��H�]Lk�7Kp��[�d����+���Z�$b�VCX<����*��Z��dq�ICJ�#��b�p���
a��W&�5��-�4�N��$5�
(Wu�5�#GB�f����U�;�h�q�ۛ������Yg��?V��E�X#s;�mu���&w��$�/E?�T��׈��UG�$�tZL���:�#ɤ�s*KCs�,�W���kK31Q�� ��6=�5�A	:;}c��a�٨P���GS�>"��08�]'�D�yˣI��a��K�T��MT����1y��EP�������^���2��߻"k�<zn�k�f�C�EШ6�	0�T�[_�P� �^n���L�[��O�L�Q��D0�fI?�|�۸����pn_~��2��_Ih�6�S�k���K����SB�q_�<�CtF536p;K�!(�)�ݓ��0T`�O|�W`/ ɶøBE)�9�p���S5{��p��~?�:���(�������3Ɔ�}�m���A�ll��%�9�S�חaڠF�8�%�����6�)x�c5ғ@(!K����-3|O���&G�y�,�[�:5f�k��m��� H
�tm�9�Q8��@�~1�nA�L/ژ-��$˕��H�0��Z&f��/Au�z���쥪b�I!Չ���5[����k2�FJ��MԠ�"-���1n�	&��Zͨ��Ǉ_VZ�z�|��<N��?�*����"}"ж(��U@�[Ż$.b���r�4�LX��7�Q)m�l^9��M��*��>/�u'풛�Hi�qmA�y���Q��Z7Ac��$fK�2<��vT�x ��ג�Z�0����<��@Z����E��c0�+�{�+�1֚����+?Eu��Ri�1�F�:Be��Yv��'��W����d����m�B2��/�_��FO@t�FzXod���xOt�)��kRlL�����S�2���5�����b#��|���SX�gn���������5/�����(�����]e�˝t�j�D�@g|�G�s�U��ఛ�'�@�D�B��a+����7K3Q2�u8.��)�G���փ`J�[���� ���+��1�E)�(*�