library verilog;
use verilog.vl_types.all;
entity alt_exc_upcore is
    generic(
        processor       : string  := "ARM";
        source          : string  := "";
        sdram_width     : integer := 32;
        sdramdqm_width  : integer := 4;
        gpio_width      : integer := 4;
        lpm_type        : string  := "alt_exc_upcore";
        req_idle        : integer := 0;
        req_first       : integer := 1;
        req_wait        : integer := 5;
        req_masterhold  : integer := 3;
        req_using       : integer := 2;
        req_again       : integer := 7
    );
    port(
        intpld          : in     vl_logic_vector(5 downto 0);
        intuart         : out    vl_logic;
        inttimer0       : out    vl_logic;
        inttimer1       : out    vl_logic;
        intcommtx       : out    vl_logic;
        intcommrx       : out    vl_logic;
        intproctimer    : out    vl_logic;
        intprocbridge   : out    vl_logic;
        debugrq         : in     vl_logic;
        debugext0       : in     vl_logic;
        debugext1       : in     vl_logic;
        debugiebrkpt    : in     vl_logic;
        debugdewpt      : in     vl_logic;
        debugextin      : in     vl_logic_vector(3 downto 0);
        debugack        : out    vl_logic;
        debugrng0       : out    vl_logic;
        debugrng1       : out    vl_logic;
        debugextout     : out    vl_logic_vector(3 downto 0);
        slavehclk       : in     vl_logic;
        slavehwrite     : in     vl_logic;
        slavehreadyi    : in     vl_logic;
        slavehselreg    : in     vl_logic;
        slavehsel       : in     vl_logic;
        slavehmastlock  : in     vl_logic;
        slavehaddr      : in     vl_logic_vector(31 downto 0);
        slavehwdata     : in     vl_logic_vector(31 downto 0);
        slavehtrans     : in     vl_logic_vector(1 downto 0);
        slavehsize      : in     vl_logic_vector(1 downto 0);
        slavehburst     : in     vl_logic_vector(2 downto 0);
        slavehreadyo    : out    vl_logic;
        slavebuserrint  : out    vl_logic;
        slavehrdata     : out    vl_logic_vector(31 downto 0);
        slavehresp      : out    vl_logic_vector(1 downto 0);
        masterhclk      : in     vl_logic;
        masterhrdata    : in     vl_logic_vector(31 downto 0);
        masterhresp     : in     vl_logic_vector(1 downto 0);
        masterhwrite    : out    vl_logic;
        masterhlock     : out    vl_logic;
        masterhbusreq   : out    vl_logic;
        masterhaddr     : out    vl_logic_vector(31 downto 0);
        masterhwdata    : out    vl_logic_vector(31 downto 0);
        masterhtrans    : out    vl_logic_vector(1 downto 0);
        masterhsize     : out    vl_logic_vector(1 downto 0);
        masterhready    : in     vl_logic;
        masterhburst    : out    vl_logic_vector(2 downto 0);
        masterhgrant    : in     vl_logic;
        lockreqdp0      : in     vl_logic;
        lockreqdp1      : in     vl_logic;
        lockgrantdp0    : out    vl_logic;
        lockgrantdp1    : out    vl_logic;
        ebiack          : in     vl_logic;
        ebiwen          : out    vl_logic;
        ebioen          : out    vl_logic;
        ebiclk          : out    vl_logic;
        ebibe           : out    vl_logic_vector(1 downto 0);
        ebicsn          : out    vl_logic_vector(3 downto 0);
        ebiaddr         : out    vl_logic_vector(24 downto 0);
        ebidq           : inout  vl_logic_vector(15 downto 0);
        uarttxd         : out    vl_logic;
        uartrtsn        : out    vl_logic;
        uartdtrn        : out    vl_logic;
        uartctsn        : in     vl_logic;
        uartdsrn        : in     vl_logic;
        uartrxd         : in     vl_logic;
        uartdcdn        : inout  vl_logic;
        uartrin         : inout  vl_logic;
        sdramclk        : out    vl_logic;
        sdramclkn       : out    vl_logic;
        sdramclke       : out    vl_logic;
        sdramwen        : out    vl_logic;
        sdramcasn       : out    vl_logic;
        sdramrasn       : out    vl_logic;
        sdramdqm        : out    vl_logic_vector;
        sdramaddr       : out    vl_logic_vector(14 downto 0);
        sdramdq         : inout  vl_logic_vector;
        sdramdqs        : inout  vl_logic_vector;
        sdramcsn        : out    vl_logic_vector(1 downto 0);
        intextpin       : in     vl_logic;
        traceclk        : out    vl_logic;
        tracesync       : out    vl_logic;
        tracepipestat   : out    vl_logic_vector(2 downto 0);
        tracepkt        : out    vl_logic_vector(15 downto 0);
        clk_ref         : in     vl_logic;
        intnmi          : in     vl_logic;
        perreset        : out    vl_logic;
        npor            : in     vl_logic;
        nreset          : inout  vl_logic;
        gpi             : in     vl_logic_vector;
        gpo             : out    vl_logic_vector
    );
end alt_exc_upcore;
