//  This file serves as a placeholder to additional logic to be added to the FPGA

module placeholder (in, out);

input [63:0] in;
output [63:0] out;

endmodule