��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&���F}���l�_���ͨ���t��-�z&���[H��M���?k��~X} �C� �6@�&�xM�\�K���<� �-�H�^�2o�k2�w/�.�S���H�7�\G����7Jα��Hu����}�@�Ɏs�����1$���CjZ��~p&qb�#
0�w.ͩ�ʢ%��lM��c���Fp9�O��.%�</�_�Q7�u�RĲw�BL,�A�Q ƶ�]OCK�|�l�}�����bt�a@��#p1i�4������I��R�T����3d���GƯ��'�����v~���y@yܷ�/?ځ����z�\WP+��枀�Wv��\��oG�e���)��!cŘ��s����U aI��hB�w�o��7�9��pb��e5}xaE�X���T]�tWY���!CJ�QEr����qx�
)irt@�K��W�� �a��ӻ��JwL�[`�;Qr��S��(���r���q���0=�d����?{Z�j-.��<0���^	p��Db%l��̇�b��A~��3�����+y�.YD���~>�ᚠ�V/�����^_?҂1�e��*~~h)�JĳF�т�x�mW��X/=� ����q��P���<��@m��]��^���'�}��U�o��-<}w���B�����Z�RX�*������k��6Sr��z<�^���K�+�(��-�wq��
8�Z�)0n2 
�>�c̟����[Y�����kl��c���p��F&�)��=v!�U�C�~և�~0 ^=�ݷu��:|�Q��P�=���>�w��Mgq&�Z����O���SO�4Hf��"�:,�� M%{v��|�mp�避L��D���p���_��uPЅ&|�x?�_6�-������#�M�:m�8�PF�����JT�[�t*3G5&B�^g�7}	"�Ɔz�5���?����cS�Ǻ��Q�A��D�&ҽ��@��R���$��B���-�?VYy��4V����0C���y�.8�1T�'��x:�x|�:+���,͜�0���U�1/Z��?μ��M`}����h�5�:����y`���4>�������k5��� �y���7��O:a9��Co}akc@�b4���sh����*5*�cȾ�@��4S��V�$��������%��So�lf8��q5
������s��_ �� �_^��&4s��G����V?т?޿ؘl�U�<H�O�c�����r�3����E�����h7����s����9neP]�B9mc��%S�BD�H�)|���WGWA��9�@2�[�Z����3F��L�1�������P��b|,-AP��&Ud?2���#ffI5ޙ�Fj��{.el���K�p/��Lh�O3��~�܏uf�����\<դ�ݍ�S��~Y_����g��TmhF�IV�(���S��ٯ=��y��{����l4׭1�?Jؤ��
��mzWq����r`[]�?\*݁��;��N}��b^�3��0Þ�i�J��8�\�����c�a0p|o�+qŢ�M�QZې�c�����Y�|ߓ��� O�R�xa3W��
�ߕ[�*mRQ�M��'%4�� ����NW�dbo�৴�V���ïg�?�L0'�?�� ]�i�{�!�lZ�����iO�� ���E$��i�%��Y����'lx%���>��z���T:��W5�o��M~�
-�� �Q�!���'b�@-�S���1,��� eP��q
.B��J�b�R?f��y�j��-��B|-W\�[Ϋç7���A�\F�N���M����[U�V�֥�]t��KLT�^)LOT�b�հ�p�	"��
�Gr��hj�^�l�r[A�ޚ2%A���9ϰ�X��<}����s��,�;ZG�����_e�ˆ'�A��_����7Q�1���X:,|�C��K2�L��"�d�6���e��q���?�L�<}�t��W���΍
aRP�k���bX����p�q��Q�N�P��z	��k�j��>؄���x��$F�|N� J�+�`|�B?���Q`�?I����?�9^��'i鷧���ؤ�G�YE�fX��1���5\^5�'�FcNq�z�����1as�Ry�k%!�f8��A�t��v���O��jgZ�40�`xt��	����ER�٧*Y��?���C;���,��͹�,�y&��!4iG}��ԓ���:�<��a4��Y����,,�L�	����0�XUF@�������@U��}�[ �d��H&L�T.�﨧�D�5�ր���]ß&KS�G��Z	���ϴ	�A���l$�
��}�y"���nT5	Ig�Y��A��<��.{&�}d���C@��rSu0�5%��"�>� �åg%�"�ulg���q����-���	�z���I~.c�ZW<H��R��ˉX��l���b�0�N�n;�J�0��0Q]bT������,��<м��[���Xt��*���a���M*���VpSh�R�J��F�<Av��_�ux�GSP� Xq�~�a�ΪB���Ry<�Ru�/[i�n8��6�|�<�QW�E@OLq{Gp�f���q��
	�.E��q����Ӕo�rM�1?��K���S�@]��ֳ�����(c���!��s���̾��6�&̠�<�zF���͹Y��.����� ��N�$�dp�J���a+��q�9XeX��4�����΢�Y�R�`�&$�FI3�4�N���I�C���e}77���r�H7�T��8P��Ac�eV����`\̻��(ڦ�
+I(� o˩�T�R2��,1Pļ3_�^8�4�@*��gb�du1#�8]�H��6�$l�ٺ� l�|���x^��m�϶4
���8�R�
�[�>s������ԕ ����w�� �
G�i���
*�����*!�S
xwkGB'���<�w�T=z���C����`�7�q�m|��L���l���1+�j>�ˆ��ꂼ=���V�ܥ�I�4�'SQ�ۓgn����a�}W���|�e���埉�������	D�3��5x����~5z�s�1Hx�"�h���手u�<�k#�7�E\1M Y���k�:c#�M�V �
��3F��Q��B��H�g�ų�)k#�����?R�7>����3��֝���-c[(�l��{�1����L�P�Z��oc͟�e��8�$P��	�.�l�7_ҡv�l�U��Qsװ!��>�vj�Kw��qu�����)^ڶ��_~��-�i�=a � ����:�x2�_ ��K36d��|��X[y>��g
�À�i�E���"�Am����C�����q�8�δ=�����&	��>T1.}�^(e����!���l���v!�.N���6��v#`�2� �f?�TJ�:-���F��껋Ք���\) �-N�&�c`��ko���7�pw���%ǩ��a
��[���粨-/�6�rh`T|�E&����dO!��^���OAq�.��8�JU��yx��z'���Jw����r��4�_ ���ʳ~���ٴ��?���vB�Z���& ���|���Wz:��u0)�oV���C�ZÅN��G�h��ϙ�3�n����g8$���L�H�\��j/��u6�����X�OL���D�?e5�r6(^�Y���x���ޥn�g�ի��ں�5%ŤQ������������ ��EFP�C���@���ǩ��7�}�e��u���)�Sq�]:WҎ���W���6l�Dɯ��ώwa���m�X֧k[�c%%OZ�� A��Og��+���V��Y�J��������0�ӏQ^s�`i��i��#�^�V���]�"g�����>)\�(�N�,s��+��""!��|�K
Aq�(���)sk!X�p�
 �G7������0f���a���~y���{_zE�Q�m1��t����ԉ�(�Y�6x�D:�#	H��u햝JX�-%��cR�qIߝO�i�6Q�D�)�"�w\��@&�ȔM�p,z�����YD���C�L���Gv뭐���uǚ`�.����o�I�����ӄn~�jJl(i�+�'M&�4�g��@�Q+�*�S�#���2B���S��?��c!L5���0�\؆�N�d��ʛ`��<���n��8��m�œ1O��&��v/ %��|��⮁*�6޳$nT?�>���2����rH�Ex��d��cH�1rs�����W50O�=L��E�|����e����U�6V���#�y�
�7Xnu���e#wYz8�D�䎿5�O_�!��Q�Q�Z�� �A2�Xޒ�B��֝8r�܇`�"�"��a9��P�SLy4>�L��>�����r�<�K��2�n����t`9��
���1�bJ跴��g�/�2T�ube�/�	�E0�i�6d�:"�	��o^�=u�Ґ����Z���-�B@��y��D��wK�k]��	�p�p훱�� ���c���<\��>1�s�U��2�d���7�\3�er��\@P��)3��041\�������#Ϧ�4{�6f��a���n�_0aR~&zC
�^[�[���2Ƅ
j6���F����9+��쯜-�/jkz4�ϣCU�WMM���=�h.�b�m���l;5����T�Ihn�n>�ųFM�;�BA����@R�x�,X-��t�|���x�rdY4*�^�������w:Njd��䍹h�ه
�}g��ٱ��J"����R����_�aY ���<m���B�+:w��ѷ����q�K$E��;���luJ��7�J���W�D�#�S���OY�
u
"�C��ɬ�-t:|CNo/���W'v�l�w�U�z��I��W�c8CXJu����$o�K>]L�2ܛ/?��y*����b�e�F��||57lۥI��z��п�(�� )�E]fT(KFK�`�{� q����uaOa��K����k�8^R��hֈÙ���2,C�p�{P��Ơi���$����C�1޾2�^�'b��V.04y�h�Ȁ����A]�}}G�
����{��zOO��Q-��&X�󟯶�_@G{�0$��b��#H`�9��:�d>ElB9��z�b�����4r��>��
r����+r~Ꚉb�r�~!{���H��%��8&�y>{ �����.P�-���,�^�4D�1��t�Q���-vԕ>���KD6�Wk�[k���'�ft���}�ꔾC`�Z��G��o�v���?@�BM*�^I�u�0wL!	t�2�4*�7~O�p�K�g�z�4xEr�Y���!�|�㚒����W��GwDuQ���8��R*+ U�,�ia�5+�y .��Y��I���ˑ@c��?ٯ0��n
~�p�	�e��@]>�(���$� 7c�KG�-N/�}�eV����]ɦc �D���_E�l��-D���͖S{�
�� !t����y:�n�9nK�]�����
���鋩��|u]g����{���ƛ�)���7�����*�u�;6~"����Dº��w�)���X�.YdOw�ܡ���9�.�!��婗n%?w_�<{zQ�M�vҥ K�'g�;W^���@�͘	���L&Y\^C1�T��6I#���:ExSm���#�m#��ŲW,�e� ڹ-�
�&gY��'�ca��)uud~7��#(B����9�P��@�χ��&MM�ްª忞/U�����09�Z%3@��	X�d�7�M�mVؒ��H=^�[_�<��h�u�T�� ���8F�Ǥ{X���� �k�H�8xdV�"H�_�����o���?e�W:���K!-�
< ���^��ڃ�q4�*"�mwˎ{�J�r��Pao"��Du��-59r�ͩ�Vg��?��D��Ș&μ�����9�6&��ۅ�ʚ��UG��$j�<�79���Z} �+!�x�2;��j�tR���5���� C�cv��e*D�^B@̓7��{?N�a�q(����֑��Й!@e�8�@Ǹo��P��<d��	��]�����9_|I�]1�AzUĩ��4�E3{!Ibגm���=zX\�!B[0�`'H�c�4�m��Oᰈ*�ć>���h� ȕEf��H�T�P_�
N�����'S,��ug޴�]���>��.��+�o���E_��?�9�ɶ$-l��/*6?<����]s L��M|0�z���@,4қF�e����$�B>/��@b3Շ��r��0<�J�k=�O���&@�w�J$0h^�x0�Q�Tٍ&����:e����Q�����Ɏ[���o|�~�ݎ�L�
�H�MBo%N�����>��=~#�v���;���Pɪ����WtB�]�b�mƦ��/}AY��m�N3z��уpv^��Ӂ0�D����OXI�ma^���X ����:��C�RȘ��%t�S�T�(1(���I��w����'��1$�M�����Q��5�W��q~�Z��o��\��5y<BH9�a���p�csD{�^�8��2l�󑀻:��0���'�;���SS���/Q��u�^/�]�Dj.�t�b�ݖ�&c���jIϠ�eO.J�.�7�/�s�!�'
�+����:������	�6��Z�<W�ʍǼb���{ٴuU[ʎ��i+A�덿&w�;����#%�����|�7UMi���M�\�`��.�Lzu��>��+���@���U��'�ou�D>�N��B-.b��ۧ͢���t��艁��(�%�x�գ3�.>��v[X���&�����I}��Җ���_r��\>��yZA�"��a�ŵ8p]�uT�0�,��~��[3͇�2��@�BMd\��9H�nf���cF�g���v0F��_�%:e�@���L�P�$�Fۊ�/g�j��>�vF��r�Ы7���%^(�fLK,��G�`Pc.�YԖS21��?}}��ht�RG��vv�0&�婯� �"��?%[�3E��t��mT}����Iɻ�+z�)�a�E`��9����3E�)Ĭ�[�LT��{r+s��7��:nFe�Hl��������K�_G��y6tu����Nz�h���7#<fU5;�/�|�ạ �\%`�oYS��e�ŭ2�!)Ù��m4.b���Mf3��/h�(F��y$�y67�D��L!͹u�Y��:��U!ȥ��+�Z��P�3)���h�)C��-nԠ݁�������0�劓V^/7j�� �)�-��)�u�����/��D�}X��7��-zߌF���G<�ع�F���-��ɬ���{�\kƿ��K<fӗ��x�qRJ}�7r��s��Ǚ<�T.�G��`R?�E~�ػ&�x��I,]���Cɽ��
��%�x����L��"C��N�w>h�
 ��4~{a��;dG�`�^X z���@a�&��v��l�����?<�˃�Q��j�S��U�b�b�L�m,<�Қ�uN[��4��p"�

��_&t����T���AY�e��	p���HZ�ݸ>�x��_��wR�4�}�#q����7�h�f ڴN�uzA&��4ب�`�u�?���v� ��[�p��;��K���H:=jw�ha���,�[��,�q���8�[��G2��;��w��a�S8�ʹ��\D�����q��R*�@��U���U^~�`��MXy��z������:��?T�s�����Ҳ ��.���+� G{u"�=|�T��B��ㇾ.@��CƧ��Gp�Z[��B��}�͆��ۃ<���f$W��":�0�� �tI�n�8���L�7������b@k��� ���bp�l-ɍ��>֧*�t����gM���֟�(}0q��đo�ٓнkx�y��Dz�c����W��Uo�Y3s9��Mn��@]�f>��tk'�D��G"�e�&��WG+�N���ٚC��`nA{Qk��{��Q!f�����=��z�tB���?��V'�O�x������[�\�/(6���9��i����ֽ�x��q��Tǽ`N#6���=1��qU���`]��-4��w뷾hX<n�oܽE�DW1Fc���)�­�G�A��b��h-R���Q���#ܹ�.�Pg��{WnUM�o'd��mE���$�W]F���D�שF1���Sd��J�z���n�k#��{�L�i*�k޺G�w_�v����a���nqe#�G�%��19�4^S-�|���2�yu�Y�"B����f�Il=�(�����*��o��$�xSU���fi��[sP�M�s���F��(���7�����Wm��\zKZ��S?��ʫ�if}��� �٦L��/5�Պ�Й�<\Ċ�z�˽�{�Kc&1�T!�
����+>����QQ�
#B��X���+%���(.[1R���!Z�������J�y���ί,��ZZ9f�xD�MA��ؗQ���:���G�7ӓ��>�9\	�]8Ϩ���L=�K�A��YL�Q([[�<�~����T�YX���@f�����}m��^l�p�n���F��E���q�Ӝ�FA�4{��w�/g�.("7l�mFZ~7\�DpW�(��@��X㼘'��q�^�&o �=����#��y�+�DRH���^Qo�{	$W��b��A���S_��	��[?��`��F_[��Qn�j�#;4���yl����� I��˹o�*�E#=V?��Ks�<�8�s��Ú ��6�R��ܣ��� ���x��<h�b�U�Uw�&&��%`�+� ��� (�@�	�֌)������-�:�4�M䂥Ѳn��<��()�_mX1IX,��F@w�(���QQ~@�#ELS6w� [W�܊g�5U������ʵ���]A�3�Ο��1x����%��m�&(��*