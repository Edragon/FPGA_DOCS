library verilog;
use verilog.vl_types.all;
entity prim_dffe is
    // This module cannot be connected to from
    // VHDL because it has unnamed ports.
end prim_dffe;
