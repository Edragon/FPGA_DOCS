library verilog;
use verilog.vl_types.all;
entity mf_stratixii_pll is
    generic(
        operation_mode  : string  := "normal";
        pll_type        : string  := "auto";
        compensate_clock: string  := "clk0";
        feedback_source : string  := "clk0";
        qualify_conf_done: string  := "off";
        test_input_comp_delay_chain_bits: integer := 0;
        test_feedback_comp_delay_chain_bits: integer := 0;
        inclk0_input_frequency: integer := 10000;
        inclk1_input_frequency: integer := 10000;
        gate_lock_signal: string  := "no";
        gate_lock_counter: integer := 1;
        valid_lock_multiplier: integer := 1;
        invalid_lock_multiplier: integer := 5;
        switch_over_type: string  := "auto";
        switch_over_on_lossclk: string  := "off";
        switch_over_on_gated_lock: string  := "off";
        switch_over_counter: integer := 1;
        enable_switch_over_counter: string  := "on";
        bandwidth       : integer := 0;
        bandwidth_type  : string  := "auto";
        down_spread     : string  := "0.0";
        spread_frequency: integer := 0;
        common_rx_tx    : string  := "off";
        rx_outclock_resource: string  := "auto";
        use_dc_coupling : string  := "false";
        clk0_output_frequency: integer := 0;
        clk0_multiply_by: integer := 1;
        clk0_divide_by  : integer := 1;
        clk0_phase_shift: string  := "0";
        clk0_duty_cycle : integer := 50;
        clk1_output_frequency: integer := 0;
        clk1_multiply_by: integer := 1;
        clk1_divide_by  : integer := 1;
        clk1_phase_shift: string  := "0";
        clk1_duty_cycle : integer := 50;
        clk2_output_frequency: integer := 0;
        clk2_multiply_by: integer := 1;
        clk2_divide_by  : integer := 1;
        clk2_phase_shift: string  := "0";
        clk2_duty_cycle : integer := 50;
        clk3_output_frequency: integer := 0;
        clk3_multiply_by: integer := 1;
        clk3_divide_by  : integer := 1;
        clk3_phase_shift: string  := "0";
        clk3_duty_cycle : integer := 50;
        clk4_output_frequency: integer := 0;
        clk4_multiply_by: integer := 1;
        clk4_divide_by  : integer := 1;
        clk4_phase_shift: string  := "0";
        clk4_duty_cycle : integer := 50;
        clk5_output_frequency: integer := 0;
        clk5_multiply_by: integer := 1;
        clk5_divide_by  : integer := 1;
        clk5_phase_shift: string  := "0";
        clk5_duty_cycle : integer := 50;
        pfd_min         : integer := 0;
        pfd_max         : integer := 0;
        vco_min         : integer := 0;
        vco_max         : integer := 0;
        vco_center      : integer := 0;
        m_initial       : integer := 1;
        m               : integer := 1;
        n               : integer := 1;
        m2              : integer := 1;
        n2              : integer := 1;
        ss              : integer := 0;
        c0_high         : integer := 1;
        c0_low          : integer := 1;
        c0_initial      : integer := 1;
        c0_mode         : string  := "bypass";
        c0_ph           : integer := 0;
        c1_high         : integer := 1;
        c1_low          : integer := 1;
        c1_initial      : integer := 1;
        c1_mode         : string  := "bypass";
        c1_ph           : integer := 0;
        c2_high         : integer := 1;
        c2_low          : integer := 1;
        c2_initial      : integer := 1;
        c2_mode         : string  := "bypass";
        c2_ph           : integer := 0;
        c3_high         : integer := 1;
        c3_low          : integer := 1;
        c3_initial      : integer := 1;
        c3_mode         : string  := "bypass";
        c3_ph           : integer := 0;
        c4_high         : integer := 1;
        c4_low          : integer := 1;
        c4_initial      : integer := 1;
        c4_mode         : string  := "bypass";
        c4_ph           : integer := 0;
        c5_high         : integer := 1;
        c5_low          : integer := 1;
        c5_initial      : integer := 1;
        c5_mode         : string  := "bypass";
        c5_ph           : integer := 0;
        m_ph            : integer := 0;
        clk0_counter    : string  := "c0";
        clk1_counter    : string  := "c1";
        clk2_counter    : string  := "c2";
        clk3_counter    : string  := "c3";
        clk4_counter    : string  := "c4";
        clk5_counter    : string  := "c5";
        c1_use_casc_in  : string  := "off";
        c2_use_casc_in  : string  := "off";
        c3_use_casc_in  : string  := "off";
        c4_use_casc_in  : string  := "off";
        c5_use_casc_in  : string  := "off";
        m_test_source   : integer := 5;
        c0_test_source  : integer := 5;
        c1_test_source  : integer := 5;
        c2_test_source  : integer := 5;
        c3_test_source  : integer := 5;
        c4_test_source  : integer := 5;
        c5_test_source  : integer := 5;
        enable0_counter : string  := "c0";
        enable1_counter : string  := "c1";
        sclkout0_phase_shift: string  := "0";
        sclkout1_phase_shift: string  := "0";
        vco_multiply_by : integer := 0;
        vco_divide_by   : integer := 0;
        charge_pump_current: integer := 0;
        loop_filter_r   : string  := "1.0";
        loop_filter_c   : integer := 1;
        pll_compensation_delay: integer := 0;
        simulation_type : string  := "functional";
        clk0_phase_shift_num: integer := 0;
        clk1_phase_shift_num: integer := 0;
        clk2_phase_shift_num: integer := 0;
        gpp_scan_chain  : integer := 174;
        primary_clock   : string  := "inclk0"
    );
    port(
        inclk           : in     vl_logic_vector(1 downto 0);
        fbin            : in     vl_logic;
        ena             : in     vl_logic;
        clkswitch       : in     vl_logic;
        areset          : in     vl_logic;
        pfdena          : in     vl_logic;
        scanclk         : in     vl_logic;
        scanread        : in     vl_logic;
        scanwrite       : in     vl_logic;
        scandata        : in     vl_logic;
        clk             : out    vl_logic_vector(5 downto 0);
        clkbad          : out    vl_logic_vector(1 downto 0);
        activeclock     : out    vl_logic;
        locked          : out    vl_logic;
        clkloss         : out    vl_logic;
        scandataout     : out    vl_logic;
        scandone        : out    vl_logic;
        enable0         : out    vl_logic;
        enable1         : out    vl_logic;
        testupout       : out    vl_logic;
        testdownout     : out    vl_logic;
        sclkout         : out    vl_logic_vector(1 downto 0)
    );
end mf_stratixii_pll;
