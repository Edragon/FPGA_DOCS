library verilog;
use verilog.vl_types.all;
entity lpm_hint_evaluation is
end lpm_hint_evaluation;
