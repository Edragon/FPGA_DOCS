��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=/�b�2uM[tڄrq��-H��K�y�L1�ڔS�����Ԟ]��:߀PW�����kF��n�A��*��ȑ"㧨��y���Zk	�Ж�F@�G�+)�Yd���Gy�<5�=��a5�1���*"}�$��(�H�d����?��iK�@m��E�9Y�[��dL`i�MR����=����1�Ǥ2k/c�<��îk�X���񭰴��e$7���U�"k.�HC�����z�� 5�n3��!�HF�}tֆ���T�3�1���ꞹ��kp&q��a�sZK�F�hfl��^g�U͜�K=Vjb>!�oy�ma��Y�s�2>N
�\X�]���3��l�c���¶�H�����R�5�6�Zi�8W}@�E�<6F\]��Ṕ:�VqW��7��E��풋.,�Hs4ó�A\�wĹM�A��w+����Oq���
"[��$�lA�-��I��=>;S�Ѣ���0�3C�|%!n�L���1�"�4���Q	�h��؞V�yu������ah��>{]��J;�]� �Se��E�eZ��\�@Iꑌ�񳕪4��,�AmW6vKDS������)�9��ֵ1ťK0&�;Q4O�:*)�$UA�Y�lT��"L�[�)b��G���o��V�������r<�k�30ĔO��^f�FX���֏�O��N0,�z��������1��.ԓ&_��f0�A:d@�p>�a��O�@i^��"��Y5
I���o-;�}eI��v&P�����V���_�1���ĝ�?�'&��{��زH� ��?�;s%O�B.Ņ0�OEM/ݱ��UL�c���
���u7߷
%����`8$0H�������n���Z�y+�n�3΄�Q�Q�v%���D�nuÅ�AY�򆧚����a �<�-3�(�I���b����$�lF�Mh�s\��B�l2���7�U.d��M�E���aɌS0,T�ћ�є�t*+k&-ѻ���8�`�Vm
��F�i�>NJ-Z��-
wI�X�|^4�����T�L�=���F��b,w	=�6����wD�A���pƕ1�r!`�4U�`�'w*j35բ�^�)f�\@�-�@zfX���&��"y�z�{GJր�r���f9'Iew�Qf���C�}��G���&���.���㰥����wQ5Mcc0k��xK��ҧ��^:Əb%��$��
���M���&���q�F&�?�H�5���� � �׌2-f�T�3[��:����خ�е"=���5)dY�l�V�eŬ���-��"���8�M;��4�lV��.[`�]i�O��6:�tvY�	/�;�pS[
[��S�?Ԭ����#&���j�1���s+�ن_7����,ٶ[�y���̆��#P ��/[��������T�n���y���k���D�%�\�e�� 5��˴��d��rYgW(&������M"�~s[O�av�W�9�(E�����˽�����kYd3����{߃Fq�%]�yK�P�O]�F���vob�#z�|�A�"1�izR!#jX\H�y�N�Ǫx�д�-{=z��� �N�5/M����M�34�.�(,\C/�ec#S��f ��=j��:���������˖K�' � dL��d���6Y�﶐�2Kp� B��[�t$��ٌ��< �AQ�����0��;�,�Kʱ�C�֤�a�@�"o�R>B�	��-�b(��Бp3 �
�׭��aE �l�;ġ��ʚq��v�,̐�m�7���!��-.b�Tp\���Rpc���� Sq����Ŝ-}��pc`�� ��h�8V�E[m�+_Eտ�י�7f�po,��(q��{N��qq�k�*Z|��f�Q}��*�X�l�U��K�ݜZ6̆��{��Fz/z-&O�����d<��pI��{�b�1`�(�v�;,q��.����9��tC�MK6�}X��,�v�ω�6�I��ft���Ũ5��P*�=`{:6��ջ8�}�cҾ�Zк��/��Ӻ�8�XiV�5a	pJS�<�t>`�.8�����:Y����)�޶�i�o��a�BrA��*d�f�d�c#�K��oY�3����/�n]�b�>�r�L�T|a`�V���j�hvl�JBc�wРCC���>�j.��ۯam2< !ߎ*��?�T��������^\���N����GcmI�n�g�~�+��	����T�m�T�d�e�օ��Hh��ʽ{��ڸ���7���an>O�j���t� f�CG �2[BD�rQ�x���#�8�#ÿ'���t�}��˿0��1 Y��2Z
��xs�OvR\�]W���`�U�&����+��29l�t�<b�rޱ�^�<!��/��߃�Y��ٞ�ֵ#L��cW�umK��H�:qt���~�C�s-�4�_DY�g\p8�@m�y'�N��Z�p��-,$q���U �n6$/3X�!ח��S��FU09(����i���Y�QmyM�˄Hfm`2�P %���(�~��T��QD�&6�kbŷ����p�Qtցk�m+9M���@x8vy೹bI�����s(��,d����s�_�Z��+���A�y'(��`�HjJ �{�j�.�y�La�3a��6/��>��!�}�y۠:Tf��'�[�*������l�hnL/�u���Mb����'�A�����;zk;��'�u,�Ғ4,���p�S�@���*o�Q�9��W�Bo���4�m2wfh�M�� �d�}Ǡ]���'g���锲w�8�*���G�c!.qGJ�A�N���W�c��7Bf���a0�߁-�K'q�%.��j%�ј)�b�H5.v`�G�_�?�,����/ڨ�]�lfix��4�FV��݂���GI���p8ys!�i@$�g�&���z3R��n�Ù9%Ɵu���/�~�W2x�`���K\�n z���j)\)T]<�~������浥�R��,U�{���u�Q�8�T�V��[��}�F�5K#�l�b!��Y ���G�е��N sֲ��(/z�L��>p����;��J.	��\��N���Z=�}�6}LA$)DA<a����� �����/�����]s?-e;nDYA��ǟ���~XgtN��U���um;��Q�qo5�q�5���o��b�T�j�8���<}�詟�x�e��S���T��Hszj�G��g0}�`�z�s��|'��4��U�>o}����}���"&J��	k��l;=�����q�u�f}/>�"��d�u�m�������U�6P�迬Q��5R����wYc������%��'<f6"7x�ߋ��o�� �����ABW��1'����^����7��g�i�s,���΅"qN�$��z��k�y���>5١t6ENco���|>��e2$a'$��jez�- ����.��˿��L��axyԀݒL$��o�\�1�'�2�F�!S��
���u��uʺ�w)�3��n 0�LxaK���r�1IP`$����J�m��n��[,E��wHd��l�]G� �?s���(���s�I�DbG\���hܙL��vK�}F]z�+9[����W�H���|�*��H������t����rJ	�*��ѯ��Cm�;I�^�����z��c�8�)��.,�4�\�e��D����4��
�D�G(�e����\�hdI�p�"��S������� �ySk�4R������o���U��@��#��۞]�]��T���ht�l)*o����oҷe����c�ZNu���T��`���I�ٻ�M{=���wiE�-6����|׷�����C��|c��/�nٷNTz"i{.��C&�*���##w7��w�溩�Z�)~0�p3"��y\o�f�r��B�����nbB�3a>-ݦ����/��f��#zr@�~/m���r����L|)Rctw�D���_T�^Y���Ά�+F*�( �`�yM'����tG�*L	9��c�iMl�"������U7����	ٶ͒y�q�n���5픫�1���<d�;W���2R�i���~ũ�u'�S�7�ar΋��*>=v��������іG�;��y�lM\�ƈ����Q�}�3����2)&B�����O���Q�U�����%b )��A?�ZoCo�y���'�H�
���bۃ�+������IC��ɍon��ӿ7 &A�i�b����A*_�Y>����/������(���U7�=</2���9I�"D�$c2?'��K<h	*�)�ni�S�x��i�W�q�UIa*k��{DH�tV7�,Y�?O�l�Q��
�[8���Bgr��TGw�Y�X��-�"T�6��I<(�����Vh�:�x��'���f~^�Ŷ�"���N/&J%��ب�S��Rw�T(*�#�5o�ۍ��R���엵�����ٖ=S""R�s4;�˅W��8�N�ߑc􇅱T�3�N1���x~0���B��ۏ�B \s|�P�XL���R��ׅ%ŧw�V;�Yj!�K8iSZ����%N��K�:ݠÓ�y�y]o��q~�_�4N���2���Rt^�s�������4�/�a�E��τ�$�ڛ����_OG��ب�t��_T���=��a3/��>�;ճ�K��~���ܚ��`lS����B�l��T���0j�u72��Z�3�F2����hA3�:k�����tl�o��b��?����)`��
f!I�C���r�]2�u(3t�p+�~|����(Ù�B4��3jȋ"��ݕ��U=D��ۄ�ɻ��d����NeZ�OC�,�e1��n;�ǐ��Z��q&|���w��h�Yt��A*?�������`�%v��'�7�)\�&%��"��?�΀�!�ʾ� X�X��!��G�H����oY�k�#%���3&ڻ�d"��ϧ�	+��%&�.}A��v�߁B\�/�VX��Z�~��0#�ZF�ܾ)G�?��aA�;BYDi6�P*3�����ȯ��J,�R����XY12Q�&�U�����V�0$X%��T5q˲޹�0�Q*f�ʠ���Y��� �X�uL�@;���ݒ *p�m��ה=�S�zxJ��xU��x;:J�f�j� ��u��I��c�� �br��O�T�|��c��QC3C�3��Y�΍�hɮ�h@�=���v9�綄;���㮨b|�N����򔕇�$�Ş)����I|�Z��W-�¸~̥	WI�2M�jNV8Oi�/p>Pℜ��ރ�N�c��rM 뀒R��p
k\���MT��fAa�`��Ҕ�/�J1T�H%�Gg0pX\m���yP��$�*��Ԇ���i͏U�pl6��H�f=Wfץ�J���w؛~�Jg�1�Ƴ��VSM�C��OPL�o��]�'$��:�n['�9n�mh���3:e_���� �ٝ�-�m��ij�!��B0\�
̩��p�cD8XڌK����W_ �`}�O��+��c+�0�5�F_މ:%3�#k�m:��u��6%����]�eu��n�B����5�,�d�tu�9B,4�7���nN:�,�����������籖.���=w{3|��g���i�ר]Ж��6��Ra�5Qt��q������zL5�&�)�$�@P6qG�(ٱ6ew�"?��F�P�0n�n�p?�l�%��%�O�"�K@�y����ӯ�O�5��ٕ��9�ǟ��,Mi�-/J�GӟS�D�/d����6�+$bq��w_%�KMCl D�F�W�=��t��A�.|���NҜ�	1��kID���ʲŞ��(�i��WbW��Dp{:F~�'J*�L�"(=�);��_����:��L�� Y�D�V[�E�����l/`�Lz�P^����Ei���¿*�L��K.�FU!�J[������ޭ��-1o�B�ALcFW�;d~����D�D�.U�q�OY(3�H���zI�[�����������FЦL�Y�M�<�Q�+(&�[�v��r�F��^~Ŗ��a����o�sL�T	��.�١���][E\�<Zt��t-�b��<�FGf��a��V��'���B�\���΄���Q��b�Y���5a=${�� ��8:ϒ�`�ج���1��I��!�ŁY�HK��cݭD �R�d�����;M��a�̸S4?]�+9ƻز�q�E�O͠m8���#l��L�'q/�ѯ�U�{	U#�բ��،��P!��IL2g%��W̅G���/{5_C�a{��R��+��ǈZ���f���J�s]��,lM[�#RE{��#�:��R�+Ab�z��iw�z�L4ǻ$���N���>�(~ɐ���oii�G�~��)3�е�ɳ�[3=� �:��B���RZ����gh�M�ЛP��zc�}���n�q�s��Tu���	�^�#�R^[n����J���U{��aJ�'7&]fr�o8�sY��c�e+�S,}�5��T�����x>���H͏�a�3�s4c���a1ӄ͗Q�Xb�8U�bx8'�J�w'D�A�#�W��S�{�U��SH嬵��U�0��3��y���<��9��<[�"A�R�Ң��`W�!ݖ�&���EcE/��/{����o[��(��E��U�0�n�O��U����B�2vR��)�^{�L��
���á�A>�X���R�S-P3[����2�<h�$v
)'���G%���f�1U�O�9�����2KK�[��'��R�!a��3{ATO��+a�a����TVu���^��, ���۲`A8S<��\�����3#1qj�c-`�%Q��H���dT��sp�at���	���O���a������2�����̛��֠��&p�#lf�o������IQ�J��	8(.���7�u}p$%�{�!v&F�ַ/��.Ԁ������{S���¾�Ћ�6�0�g6S0Mq�\]V��k77ֳ#t�]'PCJf�6��16w~��g�I|vq�.�dЍ�#.�^9Bcc���@"�'h�k	7Xf�6��[�'��/�(�>!���i8J�h�@S�d;#+	9��$������ڛ���=�z�⾾w�q#�D�8�)}��[�S~��("���Q����ئ�|�i��:WDGQjвd�����K����4� c��b�M�����(���_\8�מ��Z�����]�	r��K�H�%h�l�A&:�t'�M�W�'[9�!�%3g�@���1�Sl�v�_��2���iC���x+�F�����]����'���8���SMy�9m�B����g��`]D����b�#p�d1��S�+tA�t�@����~���)�G֚b�x���*w$>��z�ا���<Ilx�I��:7 3�e+�%Yl��*�aF:M��gm��@iuǔŴ^�00(��n�y|��iN��Հ�r4���Vy;$�����'(�#���<o�m'�QQZ��<��=�X�Ε�D�H�����b㭲)�(��V|I�T]��WΓ�լ����'$�
P��Hyz󁓄�y���ܨ��u8�Uc;j����3��)@����˾L����E��M�=a�hSd�r�ύ'Lյi�7̿_Ne+�#P`�R�N$��b�@�%z�`�VB�[+p0�E�?tz�"�j&Pv�퀕�;���RĨ>�?w�w���qL z�Dp8J�����Rပ��2����(H�QCC(6��|&�)�7jo�cۥ=1*��PHft)��,�0w4�U��=�գ�nR�$�h�|��y�B͎�DXПq���,Gy1j}�%{W<��\��|U�f�����DK}®K���#�C�3�d&��&89$x���2oV͗_�����ܶ�<�BS6���\�b���>s������D#���h��{]C�J��0Ī�s���Y�:�(#��XP�_���f�A�ğ��Mϥk�U��;\���v�D�����@�d@����4����io�Ĕ��� �T>�O�y]M�㒪IEv9Ngu��R��[����S[ns��j]~�e!sMy�<)� A���������f��Z����-��_��Ob�_��:%Gg�$r�}��}C�vxj�\�`V�yz,�:��a7SװV8s����a���ʈq�
M$��ЊvV�UN����}X�d��[���PE3W@�>�~�����Dv0���l�3��C;h9�J�.>��,��V�U_
���TM(�� �Zn� �7�o��ݽRFPOcJTeS�G�c���$��aQ��B�/����������ځ�S��"N0��qXڙ������B��F�V\��M���K�
[kl&�������yJ�g/DP���L�#G�/ƈ�k�F���=��p��\F>5Ў�P��S&��"���,��/"+n���ZB'��S�m��E.�c��jp��@;�-��.��9#�޴f�Vl��Qv���^%�>%�UA�I6&0lgqNs�3�~}��Ab��9�-*I��H��--0�c��<�v5���_���X;�eX���������X���Q!�u�4=t�P� v.���Z��cu�!O<���t9��4�U"4^�#�?�C�n����?�54w����^fAH0�xm��} ��g<��Y�� �$Z$�=��(��y��j|�d����U���j������� ��ك�Xk��ʅj�0���f*( DH��7��u�-��^0���������~����f+u"�AZyR8/bK�)�G�8����X�Y=�y8^��E_`�gY�<�m�ܷ?��l�߂<<�;v-y���E��;��AYn{D|2��c��y�!�(���V��h!`�@�%�����@Wii�^�l �9��$��w����>��\Z�"=�5;X����ܬ��)E�v�o_p�Z���!o)�$�|�'�gn~C�N��Pk^�É���/�H��=x�����k�M ]rn|՝+�#K�G?-��
�hk�����C_Ts�O�p.rs�7�0����A"�0�s���܅������U���SP��t `
ќr`2H!�����_A^�؅|c㵅�*�����SL=�=A�!k١�S���YP3^:�!b�%u�Ԗ���"�"{�e��k�+��3����@&�"�i�)�.��j\٨��j����U��>
��8� �P��>�Oj?�񙴽E�V�}��`�����|�������q)��6�Ԗߪ<d�[?�����P-���٨����OROU�o^�?�:�)$�������T�z"]��?�������� ���-��0�6Q���QR7H�2C��6�-Bq�NAw.\g�)O�6I�Z�������ԡ�䜂�s�0�>���uA�F��.=Q�X���v�k�����n	\7gh?`1�����/93֘=@�����U����0�$�W�^�̖��$�I99�=k�;�f|��(�
����G������G@i��f�� �ڒC)(�m ���V*�&1�0�7Pf
k�����Y�l��1i�'R�ɹ>���ä��{#��P�,wx�t(��e���B���m��� ��p�������l���8 �{�GJ���;��-Kd:�;w=�BSC�Zi����s`kME[��b������O'�$x�x�_H]���I�Z�#�'�{T� QE%�l����K����_��P��߽"m�w�:.�O�Ϡv8�~L�@��!Ğ�Gw�m"rl*��r��(��~N :�\�t��[<߳���f�T��^�?1��[{s�����nU�w�-��|��ӣ�n�^й�'���ȁd���^3=�0e��%{8l��)R��7`\���h�L��#B�7��[8f�+��:���.�w��V��h��cs�&���t�1��.a����	�!==[��Z�9X���Å!ƈP}(�<��]Z~%:�tPM��ʍ'��8j��;bң؂�ҟj��Z����?���	��(�R�kV�T<�ڢ�, ;�|E�1^��;|�i�>�VWcP;��Paf.��El���J5���;���2��Z갹�����f�@��vs엇�Д�c�#���x�1���z��*�|s��j*�φ�󳅎�t����|Vq:g@q�ʊ"�?�'����p-9ET����> ��2��#E�����ۢ~d�W�Ќ$q�I�����c:\֘\�B��F� ٭�U V� ��h��V��$^~�6�i�T�]�(5Y)d�~7(�3�h꣹A}2CU <���7��BҼGZ9���y?�6���bs�$��KQ+\҈32H�O*� ���s�C�~ΰ�.Β����dS�ƳFJh���M2J��i��� ��C������ɦfZJ��?����'Ȯs����z�3�����į|�)O��?��:�.�c��R6o{r�'�J�מ�贁�d�q��)��'�׻f w��(5�b�g>�����/�s2�Ć�X��
�ɨ)�ǋ��5�|�Od�<ANAc�
Sڗ������£��F��\ǳ�����T8���XQ��G~O7e`DL8�}�����;Z��
�:��X�Uk$+���B?{�rG�+��_X� ̏yc
}R�,<���v������q"��P�3�{c�:Һ�
vigVqr����x/Ɗ��R4K<CoXg��a�<����U��l����w��,����ƃG��S�����G΢TH�,O
�Yϵq�K�_���g��y@��e���y�D�6���@O,x/�%�d]�p�5��9���'X >��"�?��I���N����;<|�k ��t=>+:H���?ؗfm<�9�ƫ1��q��0��a+���
c�aha���j5�����&'E���Ӱ}{&�v!sg�B��m�ՙyR?�iu?��,�v�D�1������;�g	��P3t�ingW���� �HCb����R��5(���7�N0�8(ԕ{!�é�e?߹�hzt��3�S���K���=<$q����f��]�z��VGM���M8��� �q��L�}P�����Y�-����"Μ����p�����Q#�g���A�M��=$ց���s]�3���RW�=���?�ρ��'W@"�1�;#g�B�_�)���Yc�d�7Y'��ĳR}p_�y����Y܅6����T��ކн�2�����9�*�/�O�x]��t�QLK׷�zs���/�I��|~�A���e���my �	���,B��z����9�<�M����Æ�ǙM�;[s��3~7!����"3���~[���bM�3�]}?e4�\=h�Ug`+�w���)@��@�ռ���R]���|���E��]��c�$�xz?N�.dc����a�)��`�t���_�p�f���j��6�wQFJ�E��}�X��<�x,)�$ܦ�BBW��X9<�jŉ�$&�h��޻5��}��C1�lb����F=%���:
8	�e�ւ2�s]l�`>Ca)�T;���(9p:_0U�$�[C��_��cW~8�ڂ�׺�W0Ы}�v��0W2f�_O�AeeM]���jp�̓��'[k���Pa.v�y����6�Eu�y-B��g������/�t����I�
-�A�C�4���;01�nY��r��b�:Ni��������"�����'u�;g��6�Q>�d�~Ѷ �cl1�ooÂ�i����w�A=���ʝ8r��y�4�[Hw��;�sH���������N�l��6�l`t>� n�)�-��˳�<H$9X� �.��8����^�dj8��w��UZ���9����N���&�����E{E?���A��1MjH��;����x����~���Ƀi�����2p�)m�����R��YU>��awvw[�]j�6saA5�wC���p!"t�6��ޝ�ݦ'88w����Ow�o����{���i@�R�-[dR[�b>79˻5����
i�j� �Za��!���l�خ^P���7a"Mj���(sf
֎}�r��e�Y�r�oy�sy�ȥidw�MRZ~���7�	��Y��"�'�ܢ���E�qjql�'�/Y �4�\����`]W����/���-�tB��h쭼:;�>�^"��{ Yg`z��F��H:Y_bT������r�K�B�"��+�3���id�s��$�Fⷔ�鷤����o��g�AX�i�ͤ2�n��j>�b
X���o�<���r�^��\o�Oj���8|c�=���	��dϴ�I������Qu �˥%�{z?�
qKW�G��j����?�R��m|n�v�F�*QJ+J�.Lp�w��R0��
Z4�ʠU���a�-��&�tro�ѝ�t��V�P��S3d	_y�Þ�C7>2O$V�N��UoǶ⑨]JG(a���40F���e<"zqs��g��Rr��w(��^����E&�Q4甁�iq �$X�H�GL������w��ڠbV�Ԋ�УBaC�F�PGێ��,!�Wĝ}��Erh:p_��f�+��x��["h	��������P�QI`��ݭI���%�$�}�Ȟi�Z!~�Y��lFw�a�I�x�]lo��B���Ӱ(%X,�.��f�ԦĆ��L9�
�5Cٛ�Q�k]�uQ܎4	F�H��sd�3���!���R�d��ܤ�C��������o��X.�%�1F6�eb�I��_��"IpC#�ѻ/ò-���2����U��n�*mQ�{o�h��vݦQGW���/w\����D��Uo�?XE��/^�,��a�:={���3'�����]�͝϶L|P�H#�����7���H���b:��\^^�S�=�j@=������ӑA�B�xD������k6����۩E��/d��Q�d����7k�����O�����)�,��<�9^i�IK��A��b�L07 �k��MN���|Ŝ6�W��c_�����+�=�s����������Jӯl۹!Q
���<5G.��:G�G��DjF!�WsMҘ�5� ����2�d���@�����IZ�����<�τ6wB���/����LOuJĂ�]-^(�\
���Z��< ���#��[��BS�v��|��c��z��G�?K�;6��	s����o�bK1%N�K2�w��L�W�׉,95/�A�����̾� ]��x�qe�ї�k�-n8N�(�2�,��Z:;���a���p�O�Jߝ{�y�֮�d�|�g�3�MɐC�v�<�A���)��N"���y�J~5L%)�����W��.Q�4Ŀ�D����TAj"�*�I�/�����w����<��js�����m���(�����DI��o��'{���BOA�G���ꉕż��N���A9PWW,����mM��n���st�&O��&�]C������n�}o�Yӵ�lrś�c7ʞ�.{�ep��x1&D�Ȧ��)3a��ZS����~��w�h���h����c��h?KΝG�Lf����$0s��r6�[P�\�ᙾ��)J@�م�,t�_B�՟ཿQ'�"i:Y����|1뺵�C��ײt<g�-5� #����_�=h�)�+�Z�x탔Y�
n,�[��w��Q�}ďVM�S9Ea��#�c�\)�B�݁"l� :�(�L�7�M;C_"��л��:#C�9�����Qӛ���)!ͧ����$hB�Bֹ9�H�O�h�?���n�w�B�?��Q�����I�F%���r�o;CQ�L�p�ټ���.�O�4������Q���x�4x��_�q��r�@�l��K�;&���Ll�v��^ Rw]Ҙ>g�![i�7��^F�����-��&�R;p��A�U.e�d��٣ *o�o٪�=J ����9���o��XM���_��gf����>��F&���q��G�ρ��d�V-�N��`zT����󎺬�)-�}MI`�b��r�|����׬.�ބ'˜��nQW����G�����Z[����ڴ���1y�h���z�0u`b����X�H�a"M���@.�=�z]#��W^c�;y,��R��w@+|��K��g�0����#��?����N�XѲH�
��F7�h�,X#��y̏֡�T�R�O��z���Q�;y0���.iI"^�~��Fْq�z�1>?h�a�n�_�W�1ڤ����RB���>A'���0^��i��r����m�����.~�����G�j����!ߒ>��h��#
����\-�s�+�څrOL �J�����;�Bٜ��%�?�*hS.XXVU��r]'Z����Vd��>�6:4Ke���g.o�]�H�q�(l+$��u�2�sU>���*���|��8n�)���`迃#����b�xPզ��-W
�(�rB�>f�#��������Z����-IL�^�!�)F�.� rxK�M���1x��~�'�ϵ���nXD?���u5$�F���ȱo�u��I.̫p�	����Q�bblNI>އ���%,)ϊԻ�Yi�8�N⼖=⮨[��p�.���/%{.�ҏ��IQ�W6���J1��[����FG��������"|PU��H��B�!�g_�n���ǋ�x�F3e�gB7��^x�6CK�]r���*�}��FФ�{s�v>���vav�7Y�"F���7�a��0�b
hd& 5ppy�����_UD��o���\v'è��_%&>/�k|���o�O+�x�9AS�!r�E��<���I7*��E��S�+��u)e�Ԟ�_@�~|�~L>Ȼ�+�ۅF�Zkpe��*�B\��N�7����D�� &��q����h�)>)�g��U���8�g�'Vt�ĬJ���k�!8�|iR=6D�>�-�]	k`�"�v�n3{'��&Q'Fa�����������(����ׯ��D��Dף�ҺѲڧAk��i��à����u��i�OW���ͧ� tW��>�ZNf��N?¸w%$�ɴ��y�9��=�F����܋��0�$4�[ap[����r��A�y/9U������Жb28�t�p'S(a	W]˞������%;�x�]:�B������X���W���|����X�P���8�,	��E�;�~rK��5=���%v�����S��A%�I����'�(�t�/��Wpp95���Z&�6�-��*z�Ǣ�1m�%`r�U�j�D�X��N������rD���մ�h�>ճ��mF�����#��~���f➌�k\�&��E�Q���dx�Ϸ&�H� �3gh�6.[���l�M�m��w��Z,�L(B[]���R^�|��@��E[�T���&���-�G��	���$�5�7��#�M�߽V����W'� "���cD)��l�7۟Ð?��~��r�^�D���bK�5V��.u�F4�ݷ#��H�`|kz%\Y�[��S��c��0�rH��bi��f�e����lm���(��a�ɒP���YspƂ��[j��Ew���2K�̨=�{�})Ʊ,��Z���I))LQʀ�JRG��
ٟ�z,���Si*[u���Iam��|����|�ˎA���K�@��+h,![h������h��xF���=��A4	�MvF L#����|H9�d��ב\S�6�X�Ӊ��
I6� /4ښ�����rq���5����oH���6l(�
�*��j'f�U�8�ѫQ�^��=�s\��I��>b�'������K��dG�7��:`�f���&n�>gj����I�oF���}�ǸH�!�^ƴ�H�-�o��Dx]�6��Ab-����qO�'�V�*�z^�k�Kb�P����t�KYxe�N��=�q�^����򥏪 ���(�g�6H������\�ţ�S2w6��7l��<�3��"$���|���8��ԮI1�J��M����p��˷an��O �M'j~�(��.��7/����`���s�Y.Uo���gA��xS�>W�C��ߥ_�H˲�d��Wuρ,���X��C���i��3�w�|�V�x���b���Y+�$�YH�A����a����Q;N�f�I�1����~SʹCᇑy��w�+b�ƄY�������� �4#C��D:O�/���q�
��5��o���m�N��8�i�t�)|�g���"ꜷi8z����DUGH��F��GnT�S��:9me��T�V�Vh�C�-�	F���y�y�E���S���ԕ\�� �iu���Y={ԨPAx�;� F1��J��ܟ��!�12=�3��?����N�jؔP(R7�]�a������ҍb����+^���U��@֌)F���1��ْ/zl͔�Q�'�~;��Yv�T��΃W�b��"_�Dv�7.���������M������,�/
��!���ΊA����N��7Q���ē$��;-O���@'Ȗ?Z�=2ռ�I{��j{3b<�����^���-�I�⯎zJb&+G��u=�ң�C�o�e	�ݷc����L1���k�m??�RGCQ����I�p��(8^M��JuPAO'ڶ�sF��2r��}N��R��#�c��T+x���� �a�}���8��7 
�ۯ��w�x�e�{0���Z/�i��^&�:J�L�?��A�O�*�
3l��;eb�Ϻ\uba��W"0�l����8KZ��.���$���r���Sy����;&:DP��\�7�Z]�NU#��z��Zt�p�Z])����dm#��Da�Sw}'����"(J����ucRp�������cE��+,�␲�8�v>Q�X�eoC��ebϛ���[��zӪOQ��=�T�}��+�}cv��ޱ���엞Pt��d�\�Q����`zy��2�vf�Oޛ���7B��w�_���ٸ�8�O���B���'O�Yx���,����q�}�Tթ��iV�=L1��J�|���(8���_z�]J�AjKr�h�?Rm���#��'�
���WH���zj����l(|SH�ǒ�U�;0)�D�.���{&F�([�ԁJ�����I*�>~y��)�L"�l*��},<�qk6�+i���*�J��T�h	ѳ�sD�����T�.��gՍ:
l���Y�����sw�+�ھ�<�5r�ev��<�ۙ!W`�J\�a7
Z����D���{��y����r���5��1���>6���!�I����\kt=Jؿ���+�;!��У��	��<��K�����E��S�䲜!����<d�#�53E���00Q՝���M+�j��P{a/���N��$��5��'�͘����t
��ՠ�)$@�M��,4��`��XUW��-���#+x�
sl�O94���i_$섒b���)��A�}�����B�T��O`�!	� c�}�%Z[��B*U�=���6���Ṃex�_��1�2��m74��%?���5b7�!^2�,�� V�`��v\ȕ;��J��4ӥF�g���a��ŵ����9��dc�I�*�\�b@(��j���-6c@���h���m�F)�K��,㯟��q��\g�@�_S�����	��
� {7����d6
L~�c��Wƶ4ژK $�t8��f�C�<k�F��QH�,��*�����(xU1iк:��~��Q��<R��SS�
I �@�����|����;�������"@����K���Oz�$�!�wܲ��l8���'?AN��Ψ�@�ĥ}୷l��.&|�x���0m�$A2�="����Rv1f�<N�#���1�J��|舮=1��|d�k�V[�\�¹[�J��|25�(�KIS�8q
j+i(3�u�˗�df��u��_��dJ�m�L�]�R�V����#T�7ꞔIR�Z��A�墸	�b�z܍�9����JBls[c9PL��O��)�_	� ��� ?+�L{�{Bjy�Ԯ/ $q�e�X$��w>�X���כ�t��[ȁ�g4�í\VP^�n�n'�ʵsɶ;cgԡ �ʄXm��O$�y~�'6���t���:�](�O���d�9,:zGsR ��I���Zf��*��F�x1�����R�Ot@�,L?��o�9��l��n��b5�>)��Q��V������W�{i������V`���k��齛��u�Uq��a���vW�kE�Z�Fd��O�N�y�*�h]_W�|*Ug�YI���k.�`��m-[{�>�i�I��Xp�y��V}t˭�o�SQ	PT�NG#+�i ���$WDԠ]��m�5���;[Z5�$t��Ɯ���^:��co���Ђ��^�]���Lޮ�������Z�pb�w>�P�v��:±�鰃�c��òO�����jY���,�3ȲU�L."-U���oa, ��Ё��Ո��}˫�BQ�OB��s4cLǻt�	^]V�i��h0�9)a�{��lTF��?G�!6�04�n"F�U!�^?r�C�ut�E��m�Q�xpU zK=���'G"��B�h`�nl��O����K�a@
m%�/EmN0Q���@�K)��gt�Q�G�
��0w��$���K˯HKb��%���w흊�D"�rD2��`�� �EwC�[E�'���A�5`�	��0�7� ����	:G�P ��`!d��(5�=�J��̵�5� I{��ZYj�������W1eSL�Oss�YZ݋�U�������FN���cyWb�2/��_��tm:���f���Ɨ;�I>z8&!�q��E����c�v*���ŊȬv	��s_E��e�KK^�^��*�D�t/��C�<�w���'�7����3�p{��U;��G�!��3�݅b��؟���$DaE�v~N�{��9�����z&*�k�zv�$a�'�=At��|��X�`�%@��^+xj�l�Rq��*�3�1l�6�I�!��X�:�?7e����.�?�Q��`L�[�Qy�nu�ǫ�ﴝ�C��5�ű��Զ�+3��M"|h�&��;zM!r熈��.��G��h���-i�ۧ7@m���lS�"��=�z)����w��AB��艉V8�1�g��h�����N����'b9�(�d��w^��$�=��E%sb	������H�9�>!8��/�A:�4#����|���p*�1@5��4aB�� �c�������oڭR~	cc5����D�
`����~'�t[W��"�����'�؈"ǎ w����p��8Z�fT"b���R���ۣk;
)Sc�y_�#߽p��C-�8CY�W)�dsÅ�1=�G\1�2,d��'
����(s���U���i��t��w�.-���ZN�K����Vy�;V����	^�̛�PY� ���aR�1=N`ME]P��N�"o��V��.����&�B7܌QkW%J����c�[ˍTX���#�o�'�=�e�L�����.��/�a�������L޼.�3B{���mT�%S[����?�*�3*Ji��e'O�&�0�6���/���K�G��ևr_���l���V������"&=�$�cM�+�-�X�Y���u���k����㽮ЈT[��9^j���Hc1�@o�~O�<�9�`Tr*k�Ӛn5�"�W�}@�LG��J��U^y:�Tϭ�L���C<��@!{AI��AG)T�k�^�7.[��������O����[�#�G�c�C	���T}m�Hx�n�s���!`���ь);��nRL������:�-ͦ�����$7���?�ՀX��T�oCL9y���3c��ǹ��IJ-��ߙ�LtȉJ\0��[KuY>J���o��x�K
�Xc���1olr_�
!��!t��}n��5�mJ:gm��.��˟@��Hfb���txE̲'Χ���},����vb(-��J3o4��R.�J�gc׮ٰ->��M) ���g��!���[� Qn�M�Ѫ���ڌ�F�,6\!t	��Fe�-���Է�� ʙ^��S�>��v碞z{����[V�A������S����h���*�XȝoK�iq\덋�	q�]w����u�Č�����˒զ��/�LFp���������Þ-[���zс��v�%G�G~����b4Z��\�5#�d�竱!	���4�^��A}�ߥ��!��0�K�:6�Wk3�xt��wT	�l�E�����I���,)�2d;	y����c��F��򞧑P��_i�箏|��TX��k�Q������O9��n��T��M��7�].:���M�b�*,|Yc=�^��}[���2��7�_���6�<݁����B��t���$tź�v9�s����0��.3E�1�- I�wf>�]5���FE�Zd�����X���$���O�)��|�\��O>��NS8��Q��r{��!cXO��26��,��Z 0*��=����@�͏�H�0c+\�pִZ����P��:ù̵�}g\?U�\Pd�ߍ/Jn�	���� QI����$B�/�N��z���ؔq�� �_��h��۾SW��G�g�w6X�oI�m��Y�'�b����j�u�0x[<����j<�&>�K8�Y>��cݡL�7A���4J�:#]�
��p�i�W&A8���������\�C�� ���m���G.�����\4
�:��<�gLo!����¯�$a>:g���&�;2M��Gh��Y?�j��(��uy�K����-?�[�(��Bc�qX�t'�8#=�
]�.O�Ȱ�yU�F �c���AmA*.���ժ�/�=S��QwOz���j�[���hz�T�ÆEY���u��W�X%i�O���O��O-�z�C����z*�F��%d�i��d3�%7������%���k R�I���]�@�}c�Ũ�t�P^�Q��`����X�f�蒾:I ]�1�Y ���)�w?���#K"Ӌpd��3�O,L�-��6��Н,�sױ��@iz%ˤ�8�8��F>�Y�+�b";� _�v+}�T*՛�le|�sI)������M
6��_��0��ʶ]ͬ2�Z��"��x�qL��o��h9��/.{��{�2i9AT*�xeԦ
ḏ��_�"�<��8=��� ���������8}zG��L��O���y{C�0&-�4w�MXȑ:�L�
�#��	Lm�������݁d����h[P%av\b0Lt���}�H���!�K��y�`AzHB/Q����	4wb��.���i�&v��|-�e�*����v������K�:~�β�l����+.0@������fCc��)��o�j=װ������1����q�o�S�)$d����1��R��jF� �:�ޟo%�^1I4�Jj�"�D^��_��ٝ4ZLm��%�ǦA��B|>V2�B:xς*Λ%�_��Tk�� ]p_-\[�G[�O6x[��1��I�+��QY���$]����W���.�֎��)3���Ca_wd_c�e-\�N�-Hw���Ôa��H�,9��i]ʌDX[�'��@�nC�p6�s����+���F�;ժ�h�X����������mP�:jeE�;`l�݄�����r`[s���jEl�`������Ѩ	�������1Qw$��E!t�u=��i���	pɜ~Z{�_J�� 1�2a��������/���\$��Y��2B0V�Jq};'��7�`��9��4�94�����F�u��ҏ#P�qG���vͨ�y�g���F�m�=~b�LP�m��XP�9��G�-�1fspS��/@�uB��wGs/�j�+��R��u�ѭ"É�)�}������Д���8�oޮ��oŋi��i�$�{Ƕ^���:/�%.�H�V'�� RDG�H��d ~��6M	߾�GH� "x��RS6$��D��Kk�/!]g�.�O#�!_`<��}΍�b+
�@�^�پr���"We
 �\�j�__i�y��Bɣ	{�:`��?�������yҳ(�ɿ����-�Ug��D��T��99#� $�R��.�*�eO�5�\�-�S���!��4qT��1�9q����Q���^Rl���S�}��'B���X$��nb����Qۂ�K�Ǳe�VG��r+���S�=��� ��W�yɤ�P�+Y��/!�f[�u#�Ec��#��G�ӵO����+��+>)�aZ����x��Io �9-'.��(�Ǩ~�N����<$Mt�;�/��P5Q�4E;%�������V&=�X��'��:�]���Ž3-σ�#z��u��5��o#��/g��R��4�4�\�J�h"!I�nR�����q�$u3$�ukP�^��=2�\l��<�5��I����e�t��>�^�Q�A�U���!j���Q�_�8�s��+�e勉�����A>�w� E�[�Bk=�E��qm��Dj���FV��b�&E�%e��%=kk�[�	:r�;9�����~��s�����W{~��6}�q�E2�P
֒�II~���|~�ij��QxTyw{y�D�,��*?4��@;�aD�j��W"T���Im��|�����|Qe������N6;�T\�7��&|���!W2�`�a��!�������0�k�\ES�R�W���U^]�hJ9e)rSĴ@!��]���9h]�67F~5>
�'���>Q��G�A ��1>��Q��#���]�
����zz
(h�]XVӣA�/g�e4�v�
Z���v[e�A���6�5";�V�9���>�wM�_�{��zyK�J�B�è�ߨ�mM���4O�>�g�#8��t񖡭MBN�Y�m�z��2�;��.�p���w��h�*=H��a%�D�� G'�{gD i��+����5��ǭ[4��\�ذ�� �����C��rC\f΃��l�7������#A��!��C������%�Lg:���<0|�a��(��T���[��� }�i�^dt�Z))n3�M�K��~VL��{38�9�u�k���%LM%���>o��>q�A)�࣯��B] ߧ�b��M�tM}N�pwDg�:�B>�U��qI�@��m9o܅�Ҝ��#�������I��%�q$��k���k��=��;�m����O@����VPs9.��3Kٯ5t���[�,Gx�r�>e��xb��r��@�G[�HH����:�)�����x�	�G7"Q#~�߬K6��W?څ�:G�8��b��[�yԡ��Kh�4npWӠ�9~�O�B�恲�(�=�S���f�P�����D[�JzW��f�����OF��j�v"��uH��Z�0��lÌ7UL�}z�'Q�$���0g�6{�FV&�b���=�#W6WT�iA�ώ������H�]���A��^��E%��C���-�N�
z_��!�
hч���y��q���H�â�h>�ʐ��XJ@l�)N��H����bj�/��Z$�LG�{=������E\��L��\:�K�4�� �y[���+�sW�K���ա�����+!��v�)N��"�D�L(����M���A ������C�Bn�o��**>o�O��eM�����Fo��G��2�pD<`w�����2bS"�,v�%qu�u���E�Z���d�+�돨C�-W�u���0�(=�+	�2>��P���>C���Δ��ɐ(��TNkY�~��@[FL !g���A�[����/Q6�>������h�K��@������Y�+GI���_Qk�<� ^��0;�V�I�I�ԍ�,]�!65�1G�	|0ӯ[ ��Æ�v���z�Zw��"�|�)w*�w���3:�l2�ǁm�c�-
���t/9@K�F�
FR���C�:�zq:��r�@
�N���l+�6NCFW�ӥ)Y��^*�?bU]��G���.s�G�=#s6��� ��Ouo-�}����Kȱ��2~�>�X� �S
��P#�s@����Y{ϥ��� z�[�?2����n5{)�KO}ΨO-�<l�J�A����Q��H�!�قS��k��+h/�MI�앳�v*��]e�o�憄r�Q3�)N�wc���Ƀ�y�W5�>,���$Ѧ ��z0��}�â�͓�-jzӐt��o��}W�ChʅOBv��L2��x���5�'�DIn�^\R���	y�.�N#�'n�6��M0M�
�%;��V��5��x�2�B�������Y�s��T�)���I���%�R��R���X��{U�����0����ڊ����I�#
 ���c�C���r�r�;��r�r|�M}��㽅�2AzqvDII���h�E���`y����Q�1~�߾V^0Ҋks*	?�T
;`0�x�}�5���GKڂ��|a7�-sĐ;+�=/��Eɼ�_����(/�@G��b��>��q�+����ʶs~��هK7B��o�&�b\�@�S	N���D�s�?��(m��{�9f)�4������>C��$;�F����p�mn�zOz�V���&�iM�"F��n ;�,���N�%O�R����*���q��!��=�N���׋��D�gw8O���a*�O���`w����� *��芑dT�]� "pnE"1�<�=��.�?"ِকx���h�.���9�i�J>ihs�8�a0"�v�#���M����z�owIÜ��*Kz����:8�\年V��>q�*��g�x��+��rD�z�t$DCg��� �7$����f��3.�i;��A�����
��*5��CК̔�ٰ��%SF�9%K(a������NM�[������S��0�u��86��
�7���M1����I��%{�n��؉Х�9��l.P�ѓ�#V1<��ܡ��q$_���[@�KV�O�B"�j�=��ԃ�s/j�xݬ��@�,����n��;Fٗ|tr��.p3@�[]J�89����T���!	C�@΄�!c�,��%@^���B�s��) �����Ee2���PS���	מΧ�5�X��H�b
;\�(%U�����>P�!�F�t�0��b�8�!9��} 6�[�?6]���V���8�}�^\\�X�E�2��AZ`o�y���+��[_7�7�PR��V�\�蔄'�Z�L���
~I�%�5L���<.���V�λ�X�1�>���7��t�؅
�~L	�Yk�u�9&���|�.��?��&C�1aL���U�����2�>��/g�+�#�#���yd l+z\�Q����n"���gpx�]$�(X�ӲD�I��� ��M�P�_���-�q��
���\4	@�	���(�~ۙ�6oi4��</���f,[��	�6��)�/�yn��k����C�zI>g�P�l�5b��+^�\7W����ѬόA��i/&M��
+2�N0@p���/[o���8�.P��p�~Q.��?�y��W�Y��
*��B�N��Cp����)��E\.�Ł������2��<w����PU���@�He�&�.��85�ߘs�sˏ�-��Fa�\zm^q �Ϋ���h�4�O$�n�ïd��,zm�Bآ���W�|ҷ�ƨ�Ux���y'/��-Xcw��=��M-GJ��4�Wv����Q,4,kk�o=���ᕮ��Sԅ��b[D#R��C'Rj���c
Β�,C���8���$VC��B�����NZdg<?V� �!`I��M4$Cf6lD6zj�?1-hQ5|AV�i���9�YC�(r�H[{+�	GQ��Y1�,��US�L�DIܶ�����J���o`��λF(EoG��c�q�i޺v�V�K ����ࠍ�M��*�K�n�i׆FsG������S���-pj��[����nVN�!�&�}R��7?��+Y-P�g��z��o�Q�s�0_9��*;�����T�2��I��@v��*�9-�w<���6r4�H�ch?5��>�lGx�|�]F|����'�lqW�ȭMz}�B�9�ɥ^Ȉ�O�Ş냃��h�9��=b/~/�8%��I���_��p����zo��\�b���_W��{w'}�<���7UK���O��f}	��+���7���FTR9�V7ioK�|����eoT@ Ή[���dմ_1��>:�f�F���}�P�q���r���|Q -(Z��@��-[0�{��6s�� ���y0QG]M���f���"O�	�<Ɔ	p����!v|��o���a�\�הZ;4e֦K�+���@���+�c\���n�b�����>#�J�s* �N<��W,C�^�c�;�,b��P�\j��Z�:�Ҭ���:c�0�^�r�{�>�]�|���{j+����y��؋"��O�@y��vZ
��-bS���#�O%��^_@+�hw��X�⶚[��9�������s$u�ש �Q�w)�(�˺|����$~:�SU&��. qQ1���U�H��;��l:Z�Cꭦ�nln�4GqQ*0q�*ʄl֡;��w|���(מ���׏&�����CI�;���/�[��Ӱ��I�+��זAX��O���z�
�5
St9\g������F�O����a��xm�;,�9c)oY�s�f:��j
;���W�0��W� 7K�A�84�;�˗mт�Ui`�)���c���0R7�z7�w^s�sњ�}��Se���^�=����?�/H+�'�م=��t��Bl�nD�/�6XP�N�����D������n���SA*�#�C]�$��:Z/����������/C�t��c�N@�I��\4+��Kh�r��E�F���o|���o�j:�@<nf�`=a�͒F޼F�L�Ђ�S��J�#0k��c���2[ʇ�˛���\�.��׽L����~�K�&fU߬|�`[<�wm�Qw��4?7����p��/��
���GE��h��o/��t�*�ۗ �v��[k�ǚ7�Zɭ�Ĥ��D��g�E|�yd�:k�GjG�|!�*��Z�Y����L�s��>a`g�1�yp	�7^��AƠ餓�Z6P�⮞�Qyp"�*�~>h��I���Z���=K��)�VY�M�3q�شU7aq&�����2���iHr�Aή6��;��M�B��p��_�w�����VP��=�t0���Z��4N確�.�GD�Hk��(���aϖ0i {�y���a��uȨ�	E��)��^�U��ʤ�ҩ3'F��|'�У`�T�����L:�g"��p�l_��P���_�
2��)9H���-ɢ������l`��L�d~O՜6P�Id��X;��O�#�^�C,�g�1�Rs����q,zp0m߾�3�����wФ����P��]m�7h�x�z���
)�Q ��	�0�bf�	�,,��ћ�G��X�}��\��0��F�.<�7�2��a�j��fv��R�z������Z�'@��-C��>�� �֎��DƗh���3Dj�z0�85Z7��}D�!�V��\��۶ka��m�	������g���[٧��s�CB�a��~&X�����q:M�b��G骴��V���@����*G�����^d��Z�S=����F��rR�k�=k��ݸS�!c`O����6M�2�g���ů\����<�3��H[y�gS��R�3S���@_	��a%[�~qU�kwE}����kWB��JǌtȌ�:t�fgڟjZv�ٮ�k8��bj����|\��^|p��B��4���IS���x"�XWH���M����>©pV��&��1��fO��yX�!�[z�i�u�]�>����:|�a�������20<[\��(��k��w�Ϲ�?�o��!v�m�	�:��4�H�S�8ע��k:,&1�-�$�_��,��(G~�Z7�XƩ YfvS5�5������㜮�1�j�c��8�C׷��&��NFp��N��@��C���'`Zx>ec
�Q�Z���$��X������Ur���&��`㷲4ﺶ�N�"G��Ь����Ք����3�~��\�#˳�����"_ۇ2FE��?��+�B�����T��M ?���1��~�)w��ߐ��v��=�����]B����r-�h	̐3���\�\�-vޭ��+ &g�_�\!��]E��WI�����Ê�y���D��*l)�$xN�n�r���K1J�T�����`ھ���ɷ&�����Mn��_A�F	B �c�'Ͱ�	jAf
@s�q�V�͈���:\����S��d�v���	[� �{�6��a#_"^K���ǩ���Z9�:KF�O_5]Va�2���xLp�l��^`��f��dt�늗��N��f����!�{F��X��5�Q����t[u��pA��X3}�M�8�����C�"��`��+�#]�Mxo�Uq��s��������$=%��W!���!mA�mlȈ����L�?�u{0��Ć4V7x�&J9c����DZI�ʑ��`Ϥ�=�q�}�%�N$���jJ�?Wװv�jHj���'i�%��O�(�b)Ӽ�j��u篖u�?ژ=�Meɬa ���oH��=��R$Ѫ��_V�۷S��}�/�f�g��0���4�Ej㖞;�SsٱkN8�=��)2M���-A��>���e:eF�����2��<V�Ƅ�6�e�OD���\�'7�SҖ��N��0���; {�w�I���x�=�s��1�KC9�Z�I�TB��=�i�؞4'���Ǒ���A`f~s;�T>lz�D&�ɟ ���oG���ceW9.1k�TF��#F�c��6�-�25Eo�j<�}W6j��ٍ��?����
���L�5�����[{f�̘
�ԩ�R�9�K��,���uRӅh�Q�6�!4o''	�$~(�a%eع��ZHpw�8�!R�����p.O������1�6���@YR|��?��2����|���1Q��������x�̭���3|�����,8��0yl����-��Xg�|� rw�ə�q� E gV���Rw�A5*�c��Ģq��F�D�}�L��_��z�쪨"�U����H��(ޟ.$�`Åz�׎kus��\�_	��� dT�9=�.�k��ڤ0|�
���x~�YyT#����������$v;~'
gC���VݣBi@��9�����~,�Ƨ�H�u�%�_V7��5��)%�C[ԣ����v�x*x��N5��c�Q�M��AD w�����M)�S�l��#ٶ��}hFC+ۧJ/U!ʷ!�\��_s�1��Nf4�E�B�9����ڵh�Dp�������8=d�$��gV/��$j��ߺ@�!ߐ�T�����A�l/�%	uQ�Ɋ���:�*Ԣ�_9���|�u�fW�;܁����Xh�9(@Q�j�s�,�=�ӿ�sh��"y9����qD_I�x嶉��n�P�VP�veXR`ğ@߿� ��+��!�Nգ��&� {W�Y7x�}����[�'f���m�S�CP�Gq2�\j���2��^r��W��n�=3��R�t6�W�Z��Tq`\ć��]Tw<���f�O�~�a#"�dH9Ͱ�4w�3�����4��Di��	���Yz3;$��Wu&�+↫�)i��5�t�7 �\���.�L4G�$0M?�����n�$"��l�hG蚯�1�;��*P��e�Վy��UG��D��	�5.Q+
��a�i�Rϴ�`C��g 1te\Q��B/�M:7��X*�#���@�M+���g�V�*��[Ydu�oW�=��&���a���l+;��dcP#1��%�Sb��V��L��VU��&�j(����@3��󕅤��k�,E���RP)�z��c��(�GA"�x}{�H�����J.ۿ*j�Ρ��hƂ�~�� K���s���)kz9 '���)"n,η��/�SP�J�);��
���I�,T#S뉃|���6�� ͹�א��q@���.n���Bc.H����d_\�G`O2�M��-9�h���vQ���d�΃�n�J��wIDw�Q�aYM���#����s��=��?�~E�u���M�u���/���IrEYV����F��?`�������6��¦*,�f�6I��⍕ċ�}���+���z��� ��\{��iS5� پ�~B���^ʀ�]��w� RK��Ι<�\�¹�g��t�RA�r��8�ݨ��dh*��`?1*��p!��|<�G�J�����-ɪd����ǫ��~)��c������Vg�ۖ�Ap
�I|����;�T ���fď�Kq�S($�
� �:�(�$�h���Xс�l��P%�	xc�O}Ws���������|�m���r bg=�lќ7^�Ac�G���mr ��y��e3����=	>9�6��Ӓ��Z�����p{B��}���EK��Г��:o�����h$3��@�C��ќ�t����
?�ml%᥾��m�H���D �,��u������pM�,U��L��0��:D-�{fH$R�'m!���[��@��8J�nX"��� Ͳ�r)'b��@_��zl�m���.��x��Q8Β�F	=B�����A[m3T}���(�� �<��$���k� =[ �{ ���!.�sH��}��F t^��􂽸����	�� 65޾UC]<9�HC]кR>�4�874�o��
Jx��3��IBǣ�N"YDN
T�#���;��p
+��9w ����x!>�+&�z��be�yYN�	X.o��B�'Z��gReP��1�!��>m�6����d�ed��^Q-j��-ɢV���*m\�������)�y��Tx����ʕm�4�~�<�>�oY%��P,V@�l8�:du�.y�4l��=�q�u_�����Ak���F�r^��"$��[Ų/-,B��#�<�e�+��3M�?�� hrsx���o���,�#�[_��M���,Ц܋��*k���S�^\b�����a�W�[��k}d3J��4fΐ���4j�5����z;�-�G�����+��frY�EF�  L˅��H8��~��_O�������S�7�q�(��oF��<�C}`����u�%Zv�G{�
��@�C�mN�Ѽk� .3�l�B�f�㊦�^CPe��b�:w��W)�Lz����:G�H�¡#*�D�	j�6잁D��=0p��wuk.���0O�����j^F���\��Ⱦ�S�I S��E7F�!�f��&��^7++�H�������;���U_ ���韃��-����z���v���Ja#�a.�����8�l��6�F�}���@4oK��	���.�t�]����ޕ���,���(�FwB�3QL��8z^����o뛬��L}~޴���O"�ah������`7�_��=-�������D�'#j���������N���~Z�O�תm=MbJ�7��7o�ˬu\!>�[��k4�dXX:(w��b?1��c&��)��ϳ7~��� ����7�?P:�;8����d}�~ÿ�b��ҷ��	���=W��ϑ�x�d�	l�zL!b�'��]bx@����
�N&Q�0�6�<����	�y����2�A-��t>KNT����/' CRF%���N~\��΃�G��ζF�^����e�"��$b�~�&0Lʊ��3[͘p��D_�ǔɞtb��z�J���a��qf�d�Y!%���cqw�C�̝F�����u��7ND�k�s�/ ��C2��8s�Bc`Tte;���t�.�;ʣ�{�$-�h�E�a0��m��%+�5��l��� /+���J�*��KX��4�Zv�7����~W�R[c1�T�	��+����{I=}O�,���B��$�;L��T��1)�;�]�)Y�(4u��8�o�T ~i<%?iY�l�/�̱ �*��g?�T�>�}�LF����(8{[D�Ke� ТM�Pt��>�q��v�rSs�uD���!�kOv]$��1[�\`n-;��~�xq-�#
�?�H2[�5Y��tt�O����v5Z��y��q�ʏ��K�-u��Mz���_�/���0��kyQ��-�ގ��:O�s	�a�<(���k84@E"�oy���F�]5Z�ٙ�,.�M`��b�K�/(��dGђZ��68c����ٓ�O �}�y���./}VS���Gp1��+��${b�OkW`�{sZ�u�hА,�j�՞d���g�W�~�;�҉�s`c��S�`%R� �޽U�qIm�~�&���a�Y�~H�s����8D︿q�����%A�r7��Ŭ0ļ��_�8��?׭�U,��=�EOr��?�&��L�mj;4��(��L>PϽQ#�����d�_a�l��[��//?,_��Q#>���g�G=D5 5ڦ�����2�z�`�ٯfÇ��ᚎq���E�e]�#�7��TX/X-l���K�P
1$����n��f
�)�RsU�R���\af)�6�A=Wo�%f��Þ����/��._,���{��F���&�vNz�t�o�x|�Jɯc���B{P���J�Y� nt^K%et~̗dJo�1�{�L�q]�����d)���]��Q��o��E�r��kyF}���Y�̢U�⥡��1#bO���"<z��;�|�py:����j��!�KA]��	�n���.
����!�g���5�獵�0�ʚ7)L���`�^�D�^���a76�Y+SB�P
߈����{�*�����w$˓���A=�$���'x�k+��|2Ϊ�ǾB�TΖ�Q�8��{�"Z�V%U�{��t����-���>~��S��R�N�6F*w�A��X�Vu���P�R�ŵ�!��m�<-�[��=����6���}�f5W.�Gp`h�a���z��5��S���ykM�8�0#IF�d(�T�����U州����FM�'>�Sr�~��û����KW]�Q/t:0��b2;�%��z�Ǚ)+6,���G.�P:�.3���J��l���I�S��Ď6�!Ή�1�^:�?D0���oM�t�Ͽ��w�~�MK��{@�����H��}C�p-%�E�Q�+K��O��1+�|)���q�3��@^5��]��D���`г����'��	�v��tT,�6et(r%~^��	v�j�o�SR�#@�	�K��qv񐟣4_�B��s#�h�#��Q�3�<V����i��*s��ŴQj��~��;��l��N9"�Y>�p�G>��~w�H���Be�!�����Ѹè�Z�f��s�GS`	�DiTa)?H�	��Ȧ��u��|��î�ǩ/��!\߲B���5�tC 5/yP&�������!AV:�8�jR
í��A�Q�U��TC���5�Mu����z/��O����z��v\0+S����e�w����.~�5�ٟ$��|�x�K�T2�%��sWs\�fկ:�ݸI��H��(^�n+������б�z\�0$�9����r"8v{I�D�FZ�ty���T2�ʀh�{g��'f��s�Y�l�ԁ�|Um�
�=��-�g50,6��R�o��9M-�ǸJ�G�R�B�L{\F�a��K�ҏ�ji+�,Q�^!�����΅��QC���R*������5 x�� t��E����h����"��|�_��Lۣ֟B2���EzćZ@�9$���j�E&z���տ�t��,���E��w���np�c�Ft�K����`�)�&����R�&�DB���~��qzl�X�j�f�S�
(�/`�l�p�������7~�'�n��e������
���-�K~^r#���x2�����ƹ��J�d���"8�!�5�PY�~�΂\ȗVҪ1Uqn%�#R<��Y#p�M]������o#�j�Q�r�L�R>��e��P�$v�G��cI������co����M.�S��J-���Eo�����,���
�� ��tgj5��Ҡ�'�"곌 6\�B����(j��J��H�@�~�]��H�7$U�ٕ�J��
t�`�ƾ:��у3�;��9�5H�:T(s:��=��@�Z��	�HS�96t�{�Oq��ȌN���3�&(~��cn���g��?a�f�G�ކ�'	5��a��Z)����e�R	�Y��-�5I���j��QU�vo����P�9����S*�6��]4���s��JD�)���_Q�?x}Q7
)D�b�~HU����)AUH������'��M2߁��'͞V��`E��H�O�0D�8=#�<'�LoM�R��c���VL�w���W��ϑ�EK�[��������Ƒ�F����*E���[KŨ�!�
K��>U��A"g�A��}�$�6Nf��v2bh@ʾ,��5l�>�����n|�!}1 'D�.ܽ�P����K�Z���
��B����W*�U�חK�X)�G�wM�ȭ畑}N�3��Np5�+���e ���$�Qr�m����26�4�vR��80��u���n�~�ֹ���l|+�r�7ڝ�1�U��}* ׇ�9���T׋��Wg�6�h��g��e�z������.�>���+�\�#�t_���	�I�mE��W�mŬ��L@Y`�
[��4�6�zNʧ�"��Y�Y�t١F#�nI�)l?H;������J�ЮlhjXa�ŸnU��^j�iH�,=�om0k�r�V@T8��y��)�J�Pc��p���Y�{
$�6���kw�7�HaoDAJ�9��\\Im�!��4{cH��)��^���1G��a�k4���R[���.D|A*r3���Lw��N4"�$�+��E|~ձB׋/��I�}s�7ge����<'��_%3�j'���P����v+�ђ�	W��P"Y��c)t��5��S=�$x�]�N��u<�:�aoX��F���Bi-��p�z�%# au6��]��&��m��4P�H�d���t�`%��W0VN-�y��-$�P�o�s�28�x� ���?Tl�����T27u�e�'Q�1^��d�Յ��c��N����wjNzϑ��z�m�����[e��x�~������/��C �Q�2�̧�������5PB�Ĭ����Í�k�TR���w]<	�2���gj� ��=a�Q�K���Sf����4o{�r�����m�^P�ec�;�U���~�$�ܪH,�ޱ�ۂX6ź�0�ӛ�,�"Њ��d/#~��(!�~+5��`�6dUi�ݠG�q��ԄȨi��w|]��!֩p�7�N�s�8����*��ӡ�Ɨ�h�Wm��ed�25F���`F�
s��6�02�x~f�M�G1�(�����c�at��a��:胳��ne���h9{�@�BD�|��&m�Z�`d����n���|�>����n�C�������&��whb���^ā^�g�~�x��`k��WA�&�L�Z��Y��F������c����|foF3�%���G�6"��r��y^�o��e`Ry��,��E<s��1B��$����(ZUz�G{�l{0��c*e��Րjt�u(^��Gi��@S�_1�����'Oc����T�����b�Ѵ��b�!�4��������yDHi["�2QV��Ӱ���	b^U�YD���rk�}Yfi-W�f=��m����c
��9��ި��0!�����h�ԃ�O�)��I� ���f���Ѻ�Bh������]��	� ���
U�OI���r<�d�	�X@�Bm�5d�4O�*��$��2R�@M)�c`�:��$,�B����]���.}�t,C�`�KΣc�`e�t��U4NK��>���僌k��������>��l������l�:��q�2#�C�KE%��]9����+�Lړ�}�d�C7|Rm+j�c�m|�O��U`a�]9���2������9�-Q���l^��5��7Y`;��"]�/�h���FFa=�&le��~���iyg�T�K����
w�u�Zui�.�ï3�_��%��97J|�NQ[Q�;I��5E���)Y�����ꩍ&]Ca���S(\R8�웈'�Sm�9�5;T#�4�'�i -6;���;���R.8�E��&/[\�A�������;�}&_�L%螭ac�����џ�'��)̶ӣm%�P���n�]F�s���<�,�Bf�M����]y�x���{2Y�C��x����2�@8V�pfa@�����zg��J���Ԇ����'eX�x偏�?�$�3��
"��'\�uEZ��G�יk��'�c%�}dܴ2z���gz������y� ��
�o�	�*��C/���񁍱�yC�g*&+X�F���ͷBE�"^ Q���u�4VV��2��υ8����7�_�C������e�PU3^W�D�7鏔.��z<��C����%�	��?�D;��9�^�ɤB�o? ��z:����j�B���_��*fϞ��UƔ�8��/w?N��2�LJay��ey!q�O=���3��',�=h�! �1-�ހO�Y/�6v�e�[�Y�c����L%�i��Q���+��",-W�~�~�GdY{�Q1�(��{Z��F@칭��[%>���G�&���C���P�]�3�%t}�s�]��+�y�?�P�?]��R��X8�n����t�܅�h�:����f�y@7�	��h;�)B{H͔u:}��{؛|��^ ʝ
�E�D�I^-��f�rלe��h�18��4E�;)<�0�#!�\)g��EX�T(�ۭ)�\1v� -���횏�E�w����C�S0�B�K���L	k�y	���@�\J����4��BA>��^����7�j�#�+��A���?q��������n�t��� ���Z-Q��������o���^��v\�dЙ3ls�QMu�l0Z�$8#�`h��}��i�U6�"R�%^��#P@ߛ�DW�HIN�,�4N�4�ٗ�N�AL�[|����H��
a�0� r���nv�{���8/_����p��dH�C���c����0h��N,S��SK�뮂5?{���+|T�v�G	Z���]�D��G���Tꀣ+~1�"`7�Un��&��,���:������Td�uU?xs���Y�
�X �Odw��{O㱁���3���콝� ߪ('�e��z�;��+���?N�z
C2���W����`1K1�v}�M�,��hj\��1�_�yT�{������i|��x<Ĺn붿}�ܵ��<�6[�TqX�q��̳�����$������;WT�9r@	�f�;�=��+&�V�d�c},<�K��Q?�A7R���yH�x�nL�;|��$���mQ�F�� �T+�gő���d�`?��a���~R��2D��\�������_4�ASGfM ���x�;�ؗ�F�S�}jɃ7rt���fMf	������	y����\鎝ƀ��ϩ����;�V��Z�����L{by��Bڒ��g�)"��p���+��	[ޭ��JB�/�Ŏ�̠͍M�~�e*����k�G��+PNouo0Ӹ���ة���#ԣ���H�5�i��'5��!з�;V^r��F�
*�p�a���:�6�:HXkB?�������, ��F��_��$�r�W�(>�����k�gc�5nW�l%���^�Nc�=��[�K�8MW�{�}�W��(�ɻ�P�����q��fPi�͘�#}Զr�S���:;��4N��^0�yY!FFkl�D�5�s4Mۖ΁��_D���a���eCwNP�tR�r�s-a,; xO��&�Z�M]/�*�=��?���3���ym��:��0^R�d:*a�������:]��gM�G�Sč�XPz�#
�;��=�?˯OS��'1Fd���b9�5[�������Ǝ���Q[N�z�w����nԮ��v�Ue����Z;>Q4O�t�=ڀ�3��_�Ƒ�6�*<,D���� ��1��Us��1."�C$�0�#���'@2�bq��w$�nU�ogG�}�v�Y�DO����݁��=��,)�U0c�����BS$�g�^��6��{�`�;s�d>&�����g*��*E�~���w
'�ԗ����z��V*(g	�}U�a�Y��$��p$��f�e�Cs�M�v��(�<�3o�N����ň�Ov��_����7Q�i+eO���UNd�<�ZUo>��*�Pf����dY14]�(���_o[�:ω*{!�\�o`m�Ȉ�&��s�X�Γ?��?�;�~��L��q<y�m��i��N�����_�4DT䯁��P��9��CE��Ch��'L�[i������$	�Բe�Ց�3=�fl 97��R���H�w�!�0�n���}g,���ORZ�iX57֤��*2�64= >N��|�=�wڟ�'oL~������ ��iS9����ZC.��E��Ve�������H�`��?�i�ռe�"'}Ff�L�'�[�J<É0��r/ⶊ*���Q�b��q$	L�5`h,b*h����������>������q�M��{Lt\���Ty{�H��� �d|_��B��E�z�PXT.�4T=�59
�|1˥F�Z�P����C3[�d�)�/�3V�ӧ�#�G��ܐ���QeRA�Kζ���]�VQ�+���br�f-� ���t�WxQ�t�N�,�����|�H�&��v�^� dX��+���m�'j����jI,u���Wg��e6L-N�t)(|!�����?BŋYAҨ��B�Zֺv~	Fm]Hٞ(|�tuHg������O�"N�܄�?S�i8��u�e(R|��e��@g�n��@��b=-}�k�T~�cY �>���j�#:)��O]�~^ɘ<�"�vr&��2�y���oAC�b����K���2�<<��L[&�ƥ��/��R��� ���5w��a�K6�욨�)pL�-6���s�ů��X��=O�lCI*}1_�[�G._n��(�?4�b��@�0�E?��%z��3W�;��H� ʱA�.���5C�bs�c����tG��UO5wVot���W-�����{�a����D�~A|��ucvt�l$D����3T-|�-Wcm���:�N\G�6l�I�Xb��x�ч��9��}W���L�}P�+���2�5!�!c'��Q�Nw��8 j6�UV����fY\�Y�k$�u� w��N�dn��xu��{ϝ�}.(��9�Fq7�&�ü����uh� �Bh4���p�g	�vl��
(��t�io��x-��P��w�� +�z\�a���8k4�ϡ�����Ϊ��SӪ��;��v����7X7.�U*m=�b͎�́K�)r���M{�k^Ђ8��R��}������H1��҄!ZY�]�C}�դ�����X0�f��C��k����&{���Նt�7����5��OZL*q�h�_��Ūa}�)�[c��>�i�9����ZI�i~� ~��{⯱E��;c��Ph�]ʿ	C����j-�93ġ ���s��K�zĝQ�2��F��Hkuƹ����g9���N;�l��Ŭ���n���=H���臐���{o�t�v`~��=s ϩd �� ��$���x3H1���Ss��PwP����@�1����(���N:G;��N�]�v��[r��h�Ͽ�r�8��A�dߩ	
F}Z���.FTșt��<�A��a!Zٞ����#Pg[ni �����(H�R�!���ͧ����c$V�ώ̊% 7��$,ƾ��V���~q��0���e�F���0�J�Z��U5�3����6w���j��"����~@��x0�����G��<��I�T��H>���)=E^��gw��2��G��#���xM� �n�5��Eg�q�ϑ'�/�}�XN�g��-���BM�&"�XY[�xg�]�ginu�[��wxYջ:�}=������nmȱa�ۄ��O� ����-�^b��ض��{���lF�}W�����DnX�A����u�N؁��o�k����B���q*U@J���U��A�=!�s�n֌q�R6�=��F�c_=����>���e�4�![�q.�IFg��.���|�ޡ�9����K�� �QnO�q��H�gIT҃ ?��YM�Q_z�P
�`Ȯ e����6��H����Z�T��$Kp�=5����X��&�pG�0|�j��G��Oj�K:� I��R�?B)LiG�X��ڵ�%���b��Ǣ�N�4��@���{�ΰ�oG&���Ee��:#M(�'*�Q����?itE��O�p-N9����cE�}���#�󬨾+	�LڻIZ/%�}V �Sɪ��p)~�J\.��/�J����	�q��>��L�"�l��[���`��KH�����7j�DYc�t��0���g��z"V(Ex�ʓ!�52jEl3�_'5�t�Y���>%�*�
�r+Zt���JѬY��0���8M(� �N-�+�܃���rg'"��x���Ք����&+('�?n��ݙh���O�Q�E^��I?�,�����4�������J���-jE_q�_J������V��R�c<'�V�
�_�i�6���_��Dt�k}2��鹭�Q�$B�Ό���Ϥ�jo�P�k_Q�{��*~/Jd��ϻ&'$�ńqSYE�mJ���pM(|�ocwNڇI�D�?��ǐ l��"׹��d����b�O��r#�NA��	�_o2����Y�IM{�F��'��E����s�A�dT��.".��A0�+<�)k�L���{g�����S?,X�k�7l��4��ݣF⦱�0��5�_�Yli�rm8��A|�ߕs�Y�k8���m��#����=KQ��#[~�9�>� .A�?Pn�d��L�����_�
�X��Ly��9�Qr̓����䪽�i^V��]�Hw9n���ד�QD���	<�ǝ�&"4K�����B�e�Ή�?�NӲx!ߔ�>��Ȓ���h.�%��ݫ�xy�)RE?a�/�3�苂�ɠP�&�f�T��*2��r��(;���Z��?i�a�f��U0A�_�Z�]մ�m�c'bRs�KO�7�ўg��f�%hK>o�r����&s�A�/���$�c. ���{�����`t��F��L�}e�M��%�9`��4���M��F(���Őh|�Lח��Oe(d���p�h06g��yvLs�~gb��n�?4/B���?�g���0����[�'���z$}�B�l�J����Q�����ZD��x�_WWR4^{3
�{��JA|�-���R�Yc��9��W�j��FSAD����졕�^1S��j�d�7��M�����ꗼ��<��kY�t'�Hչ����a��ܦ�����7XK��B�C,`�:,��xj��*����Sc�9�ǔ��a�ϗ�'��?��+��,��Ň�P۳*�g��1��,�u�B�^z�Bj�]*%8-�t�&v��"}QZ��9ec��E=�3 �^ZJ��u]:}�o� �̓�X���pF�[��Z]59�}W�硿�ҙ��6�!o��%��y3zU���h���Q ��ߤ�5N�Cn���P$����T0�3��X^%�H~��������ƀ@�Fr�'{v�����:��CJ�6j�R�Ԯ^zV͌^߮D��%0o����I���ZR{M��!tG��A�T�A�^-R��C��4f'f��&�r�=��|�]#���N��B��<�����<�e/�2 0�N�O�l��8�|��[(l�$r/V/��r��o{kTS�����C����覹Mn�l=��Fr�{������˙b=�1��FV�k+Ԗ%�j4W��Xnכ���%�Q�l�4�[Ms�a�n�WZs�	_��pˮ�F8���˴� ��t�?�WR���#�N����xB��G��;�RF!c͑���eyKQ�-�Pev7D�4C�����SҥȚrܴ+Ĵ`�}g'��3$VM,,f�!\��hx��|r�9�^�F�H:$N�n��)i\Ǿ�I���|j`�|VA9�tv������3H�b�Qp�=\P�a�xS���"�7l�x�]\�����>��>�l���?B�d����q��sD�[B:�$�|�v�cxef��8?��4iց��}��צqVEp+;h�����C'��	C�U�4v������8`
T���4���9�r��=�!��*B�����7��[�`O4�5�=?���Z
ZT����/R�Ɏ�`h�(�����hc�2������e��N$�2���N��cʮ4ja���>,�%�"��.�&���ZT,��]1Al�$�S�Z��i"m�m�T�yVuF�^A6޷�q'V�Io<WJ����uQ��p���gr��-��-3ɾ5��h2�\����A���=WR>�~1�`ޔ�CJ�kU�P����@��,�&(����uwj<0�*�F2e��K4G�dl��Y�P�I	f�,�]Q�5O�b�|�\`�a`�����D4����l���U��P������(�c,��]��ge���왬}z��P`�/��`���a�5��9+jY���d�$0Eg�I���'�!8��vP<�9��wU*�/��d�C�y���
��'��}��6*v	Z��j��H���;~
�������zXY�q8�K���k���-��%�N1;��2��]9��ѫ����ب���U��W�.%�I�����1�^��'ϒ�o�/���4%�������z�l�Lt��~9Pl]�Nf���/�׻�x=hs'�� :�j� =N{XLẢ��05m���ٔd�EO2F t�P"@]��Av�
B��1~4O}�L�`��+vw�>��WO_@J�NP�����,�{�"����hV���%��-;��z�'e��g�����j��n���x�,=ΛY�;�:
}g�o3���dQ�����Q�ި�c�Ӹp� �P7���Xj��n��F�A�Ӊ� 1�����d��@Z���G.g�dLu�&��M�����Q���.GF�yA;z���Ŵt�(�?���-���)��,LS�X����;��7K�Hh� �$�+"�#4�j�ɾ9)�����J���wh'H.t��j��yz��9hf� ��0���]�SH0��i,4�ps�~��c��ŠV��4��:X�#�Y`y�S�w]M�J4/K��E���砜�l�T�0P��c�����1�?�2��U+�=�c��TF���,2����/5��t@�`¢_����Z&��]@�M��R@.~��≮�b긆?�B0 N:�>xZ�Q~���j}c_Ff!�0]�.�������N���J��j�օ�8�͑f_���o5s =O�I��n���0r3:<��+	=K ��1����F_��Էu��.��Qb�Rs~S"p꽬a�"1�������xGԡ�r������: �Y	�lTR�6�oS������oY
kGS{�\��;є@���Z/ܙ�%�K�3����'��V�в�:nSl�� =�Jŧ��/B<N��9��#��TF�*a����Df��	���J��Y��kY��������kc�Oy^W�:ֻ��
mBZ)�R��se��P�j�Q��Ѕ��H��J4�3���zu�|��W�\�<��|;���Dc��<Ո��v��9nm��(�=4s�އ+]�a>"�g$-�m�b�5��E�U�z�8Yb�%�˳_Ճw"
"���:�Yg�%i����.�4�h]V��ٕ� -7={UZ����n�G�������Xc���xu0f�ZR�.�ս���b����*;������B&�C�(�[oZ�����J��!8�N�e�)���M��m��M᧧o��qԪyEѰ-�LIf����G�$9�Q�gڰ]��q���TQ3c� ����G�S��9�|���	Y^�=X�{�ڲSj���}����C_���4qr�Jʹ%̖�b�q �A[b����BI]�93��Zȏ��sp!�A �ugf��i�TG���7�>�%��
�1�]�3Sw�X�t�q� �/�5p�K��gl���1@h�|ʣt�:_*l:���Puu��A����Pç� �T�؎s��)5f�4"���\��{?L�&���:Jߦ���F1Z�|�Uj"�!_11�]~.W���IX#��-�����h�xX�O��n��>ǀ!�Ψ9�m��Nz$����=4�����B�M+�����~��?��;�Ȯ#!G�X�;�������~_/qL޴�mW#6wы��\�����b 7p:���j�;�����%A!��ν+�V�2�'��N��ޗ,��H�I�I��j� /5HDo�y�w7R���&y@p�a�W�R���o{�+m��x�bR��������k���[x+� �{��9�8!~�X���;3^��"w>�� T�J�J�?���uc�xw'���ֺ��R�5f��=7@���zd{�*��=!4f�2�W����K=w�a�1����D�<�&u=v���E(&���5�D|Ȁ�X�!�ޗ�k�A�[ۯmE�対���Cp�Z�}�ltX=-.m��C�<)��}�B�@秫O�Qu�#��4mT�U�uOI�d1%�`�@*
IY�Q�nL@�?,���j��ϒYY82��~�V7&ո��M��t��Vt�YG�֙)��t���n�����/���Y��B�5VoN��I��Ԙ��l������ %�F_b���������cN�nt�TǼMbo�t��fJ�?z��M�{�T;�j���tGC;��=N$Ҙ"/w.�ˣ�JC�I���������2��M�~����y��kᕩ��GAE�b�sY�B�������&j�-L���	�[�B�Xx��9�u�Qڄ�G��ey�5�&�l���$bp[��QXn�D�����"yM@�V1����<��^�����x7��zڥ������٤��i�9��r�!ƥ�X_�1ʇ�W��R�Ux'�0��S�RO� �#��W�&?w?�'f�>��F}pM�?�Яc�!�^�E_zK yMv����.����gY�m������J��в]cB.��f�g�CV@�Ic�����]vҺ"��ap�m �b.�7f�-djIt=�~!��J&�v�
~w�~C�q��;��.�4�ެ@�$3�����2�H���S�Ԩ=��c-Ty����U��\���8� ��p���U2 C%W��g�����=�=_9( �����ovD,v_ ��#���̏����a�@��HC��>�3{�^����#{S��=�΄VVcM��ٰ�f���Ŷ���.� n��/V>��AALJVnR�������S%�%!�[S���ϳ�p0*[���f"yݕcM�:V�<ČB�u%0+`����D;�G�Ok�<��ړ�@��B�[��/���y�g��~���5�ƥ�
�;r��5���@33{��̀�C�b:Yz����o� c�:|K�j|6tW|e�(ԳPP��\e��TAX�"[��N4�߮X��?�ZrD>�`�s�"FY��62�k2[�?�=/�ض��w�ØϿ���0Ml�������a)��ɀ�(�f���K�����1�l��<����~Ș�'�����_g��:\�敏�Ф2yd���z�V_z4�^��ʝA�k���e��?!v�h.t� 3Td��t�m Z���0�� M�@���x�GJ�\�KW��B���Hh�ތ��ݥB���^�t�6�Y��O|��مaP���Dv�� �yp��W6O�9O&P^�5���Jɂh�����BS{N(���GY�׊����kB�qbj�pޡ-g%1�h��v,���Hc/r���I�!�+?ws�y(�{w��pM�&C��v�0�B3Wͅ�|l�cN(��-��Ӕ���U�;�)I��������oi��H�M>-�ұa0�SS�8�t�k8�����6:Ⱞx&^a\���WY� Q�A����ljn�N�<n>�mJ D:
�~>l�Õ�F	V�V{���$�`�
?���O3�Sa��$� ��A}��S��Eǩ��\X�25\f&�D�� 8�t�|�~V������j3=�bv�cP<��k���y��I�K�:�X��mXA�>�d�q:�;8�q�����zpII6
6v9�NM����+��xߏ��_�6d����'rg� ��]�w��(��'oVY�"�xYe�U�Y*�j�"�wC�%��Q�K����1�<�8�̹K��$jy�󳊾{��,�f�M�FիsӾ5�ѥA�jFx^
7`^~*r���Y<	�#������wb4�
śt������m�K`���m̳�L��7�k���e-�5��6�_Е�V
=A��RA�}&?�ZCi��:,AH�������K�XXQ�.���	�Q��.o��4��Z�^�p/Q2b'H/��h�\&א�lv3�F0�����ƺ�����G���C@�L�0�L0��Պ=z��i`Y��ߎs��#��h�;�p���:I�4�*�_��&W�n��}����4N�"@����g��/QГ!_\�a}HB���v�|Yg4�Pإ��R��9�`GY�䇝�.'�B5�*��T�B�_Q%�ز�=P��� /_��y�['����!W DZԠf��CY����Rg�p�7e�^g����zL��XW��y��\��>t=�� ��g����uT�A��9	���+�����5��u�݇�}����=�IG�߂�0��bHY�#ϟDR��Ul���P��*�@��o�D�\�e򕴵8�KK ���n�e8)m1�y�rKg�� ��sw/�}�"����L�v����Z���/o�m�l��A�
B��>�^�8�$sC�y��?Q��獒�5��Əэ�MHG�I%2��+1°'�TcIo�F���g��"ݨ��1,:�(����"q��(m�<���ۅ̩�W��i16���y���O� ^|�T��:����r �!l*Gs��EwB�_�:-�G�L����C;���NUbS������ߤ6ǰ�;M�|U�6ة��(�6�����tZaƁ��t8���@�FKJ� Z%�_�ތ�2���M<���`��uO��N�����j�8���8����bV��K����?�iX����!��`���\4C�b{�/9n�y�8X�i��ӈ�"���vQg�	�����=�ܠ&���"�G�uU�?�usGȧv�����[�"E���C��+��Q�\ۄ�����-�C�Df1=>ucǼ��EDC���W3��� ,E�[���z��O���ֈ2�Jsk{�)$�d��������0��>�5�h��������+����	�ʞgA��
H�<�&�(1��֠��ZN��(o��$,�YSp/�K�%�ʻ��TP���՛(�I���\���WJ��a��t�b	H�S^�R	��Ʒ�}�f������XU�A6zX�|��h�&f�]��u_0��T�	!�Uw6��
�$���)3qU`ә;Ta[��,��kWlk)_c�59̀	���z(�B��.*`�$�_�Sa#!�bo��E1�_�65H���0ū�9�`�$c����Ϧ���%p��K��g���vc�i�q����@m�:��������N�:uHF�u.J2���rN�0�:$�Q�H��WbpYo���ˆ г]��$�g=�Gx�8�(;��� ���Xf �̝3�
W��#��h� _ ��M��8$�-ӵ����$��`؝fX����|�PM	d��̿|�Iº$�Z٫���� �ܩ�y��j-d���6|iC��
p�K�ao�� 	v���9IvF/[�*$L�O�XHX�Ev,��~�"�f����(w'�f�)�"]4�`�/!
۱����J�ň8Ĺn�	�����)? u�����H����$����㝊\'��4������gx��
P̧!O��\�D@���D�j.�UNt���]�B�M`�W >N��S掷R�|̵ã�����Su�4�b�mm�M��F_1;��Jn���	� ���(2Q�?h}p��u=EOQ����o��6׀��q�D��<�&�}kF�o�`(��ή�̜�_��d8�f�jV��k�,k�#���9nA���[�Q�͒H�&�������]�`�
��F?��yn�@��!()�3\����#YM�������֎�����]��Wy��mR�,'��^=�Q 1}���"ҚhAh���=�{��-����X;QX}Ƃ�-����.pV��5�~;����M��)��-��(=�T����uy�ȷ	�(�V*�|����w��|&�"h�	|D��,*�����'K��լ�(I�B9���/�d��ʣq��(����"��x�p{!�i,P�Z;���Mg���vh�^��5�QtЃ0�����>}�$�7{j]��,�I:��їב��<�C`q��pϨ�����v����X�|�ݫq>Rs�3<�s�B���N)����G`�ip�!ډ�6n��貮!�F���t9�rZa(, }ۺ��"�W�����NL�5Y5����R��Aנ���6�})q4<_[|/չ5�F�oT���?�������کD#���&/�#��D�)�A��`+��l3_���?��o��F�@��n@=�P/�b�d ��J,���AC�?�[�}�
ԍ902��i9 ��\k�Xj=}����tpG�ݖ߳��%�c�&U�����e#ϡ'��7��_�ux�(�,��|2�5�ki����oU�I���2�pR�*����Q$��JR��И�
a8�2LѫgJz�#��+P�M��M��M.)�o6"�Z���\k��b�M-�6�C�b����~�?go�9�q�(�g�����6�tz k..q�=��d�l���!",��؏42Kw�J9��Z�.�����)���a���nPe�1?G�Ɠ{p�~9�?)����{cc]��쑕ms�/0�@Rqd�wT2'3�]����'{}��Qc���V^99���(Z!�ą��:N���|����1��n/P�����Z�k?�I[`��~"��"ecZ�?��1��$�;/�� I��K$��OJ%uO
_z�eo��/��xC�5#E�<��M���c(�7@i�F�E^پ���"Qp�h�OI��EZ�T���ݴz�m�2�:�QX���C�v=X��mX�g1a��^A������O�j޷�S6��%������E}��	�$4ލ��ÏT���s����Q��j.��w���U�ƃ"Z~쨣0�&��<P�_-}�vPw�"���������zg�g�G�iw���!���.&)2�3�$nE�_X3�ຕ�=�rW,�h�����1]��d�Ș��~�/*��HY&�pg6�x�Ê��Gŷآi\UB3�"�y^�QX�=e8SD�BM���K�KQa����mu�H��Z;��t@�6Q��v��3!LG�OS�q�|�b��U���צq�a�ڋ�%��`�SU(�(,�Q�o�Fq��?�F�h�BSY' np�d�_���P�=��䨠,��$x�S
V��_�F��g��ڀ��i���[���㔰 (�:�$5s��F��v�9ެ��t�������Sݙ��Z�Ҋh����`@��`�Ž@�j�����ᮬp�Tm���[�Յ[�Ō�O"J,���E��G�o$�Å��OT(���H��7^�x	���=�4��xhz>/ �9�3� Xkz�jo�XJhwR�㈽��g��;!F�6"�)���<��1�~g��T�4t ���o�b�J��ﭫ�Qj(XN��j]���گ�c����e|H	$�/xy�䞓~5��H|� �@��o,N����^�Y��nfy��­ͪI��aM�);ֻ~p57#%��k�	V�3;��RJ��+��*Y�>&���A�a����\��u+�l�c�Ô~���T���.+'%��N�:|eɋ-	C6ʩ����jWq�p�����WTq(H�W��X@U��
�����:ˋ����P=����8S�`C��¦F�J]<�����]S(�a�^�=,	��'1*v��q��o~�ɿ��%)�eA6n� �n{f8�oDJ9�E�J�0 )�x�o�}�Ex�R���b��*۬5��"t"�֑�| ��nւi]ux68���T��d��,��\/�a���n�e����ݘ0f��G� dҡ ��� ٓ��߂��Fu~��&dq>e,��.ᆟ�<n���ʋ��r���$]ە��l��,���/�Q*� T����Q�@���N��b�Bf
�z��:pQ{^� ���v��v��T+ݣ�����a�q�jnvZ.ٲ�,J��T���B6�����?}��ߚ��E�Oο��r���0�;�\�b����(�c���(�@(��vu�=�^+o[�f1̞T4�N����������d��]����tuP��ٔ&����]b�ǆ���ԮH+���o��D��ൾ��cq��=��y�������{
A�r*��OD���QI�`�,h XQ�Ӫh�.�^�^""2��I���޿�s��{)�<�
���XR�4���C���W\a�o-�^��9X�y�>N��{J����h���ϓ?SȮ0�!{��5Va�\h�_{�-��>V��u�G}.�!��T#�y�@�� �I`��{C9�@��}14�H�����5�cpzlV ����g��z�?J��
"ϳ�|S���
���|1b��G�&����a�;�����җ���Z�����y�X�3�yKk����_��N�L�V�-��;9ּ����m@	O�������)�[����%^-� Ʊ
�59����х��*-�g`c���\09&c(:	�ֹ����?�5� ݏ������������ⴜ�40j�U�M"u�q��"�9�N��0p+!4�3EЏ�~��v�	(m�ɭM�i��G�|d!);/��6���*-�it��m3�%�}!���>�{΅y �) ��ɻ&�!ɬ�#�V�3K5���cz�֊�_�i��|�k�Kq��"80�+Zb27���)i�ƽ��W�q��c6`O��,~�mSX�@ؤ1����*?�G��P~�i.��`C	S.��i gL3���P������2��`�x_>1cw�V`xuGG���^�	�1��AsQ��zBˑc�F�����������Ӈ����V�]�^��Y� �,[7��ٓ��	X�lhjɖ8���v@���Ţ�g��&��6K�q�}	ɚ-�l-�|7�J�wD@v�]�^���
���r<e����"_�F�qvP��xv2Z��4n���z�]�(ٛB8ԚL��i�X�ꭔ0|]&J^��5�h��: ն�d�+�Ļ�kz"�� #\��!-��GT���E/N{<�/5��Zs!m��ݻ�O�U�}+�������{%(���I㝁�<Km z��<�;�i0s����d��;�{�`�_�f�N�n�!�W'��-��NX�)�:�*�^y�s�v�_�r�I�XU<��j��4!y�[�@�cɧ��j��=4s���5?���=-���'�06��Z�I]&�co ��*;�Z_��Ek�ah�Զ�3�{�	�ֿ|`�)p�w=XBl�Ɍ��ɧX:'2[ƁW��솚pAR暖�iè�7 �jw'�4��ؽ�eyB��a��j��b�	�\����S�}3����4J�L	��� ��wCf�M�gʄ�d�X*_ ��?I$��e�������w����K�(!bs�l���_,@p���(Nf�g��Lt#�Y��)9��-*Hdr����0���d&������*�aʀ��X�ۘ�'r�?6W��)PF�*�,�r�8::��K�9��nyLluu�b�ǆ�Zd�x(�&$�N3ʱ�5 �2MI����<a�vd$�|���ȑr�GS�q�������&t�o�-�5x��k81Lw{�ֵ��o]�$�z�Ԅ9l�!��t�����Ѻ658���ž%��>M�Ep��(���W��L-�o��_A����w]l�+��*�&��A���puG�u��VpR�X��tu*���/.�^IӒX�bÞ�ǈ��K�����.��4�����G�*R'}1�ij�I�������/��qubil���\�
j��p��_�T6x��[p˖=��Sڰ��K�|oN�����/Rhz�7��b��%Mq亊�s�^�}	4��h�r�f�FݽI�f��Q��Rk�Q�A�ZTH��"�Յ�3�k���$�,���<�*tx�@n�ńX6���G�E����9{��Q��� L"'�}�i�M��֪z�L)��f� ��?��R��XZ�_Y���HRL�(������n��)]G+�],)Z�!�IJ2��J�H�1d9�����>e�IO�g��̠��l����0�9�T�0"��<�����̞���R0���ӧ����f�~2;�Z�̏���A�,#U�w�O����7���r�X�0��D��?�c�W`|���:߸�����np���Yn��T����>�U������߅6���F�\�);�kC���	�
 ����4�����噸���>�>K�5�m���HF8�>(Lf�4|P�5?
^�F��pH���T10TMŨ�����q��
	S�*��a��ICgp�i� � �w�P�|oz
B���v33�v�9�A-*wux.��C����t���=8J�U~Ê�6:":<����fF9΍�v���G�dw^��{_��v$�6ɐF^���%(���-m(b��WS�P�4#e{�j&�`1g��,ߜ�=�J�F�s�s��q�g)�s*�I|Z�N���X18��JE�q�z �ޟ�����K�`�w�JI�Ⱦ��. �Ԝ�|�G4k�ô27���߄WͺnQ���+9�0�w8�&��sгH6��h'd.���� �B� ���=�l����RZ��\5������ٹ2�K�=Z��';��[���d�X:E^�ލ�x��LÉd�E��ޡ���2+�CVk���-C�yH�A*�c/$H-�y�U��JE��d#pQM����\���£Fz�^9ڹT�p�q��s�i�M��O�xm�i���~����a4*F�4�i���xI��*�t��z�ˆ:F@����i�'ϯ�˕g^��1��3�D��-� �DNl{��{v�W0����d["��(�����Ⱦ5UM]�iR������D"���-:J�u�,I��D�owH��. |�J�k%pJO������gT���1�`{c*�2<��e!�{- �\ �ȠyX�����6�lBӶ�Fi���a_жe��-�=�N�*/�e�k.t���+�U�-V���/<�{�t�j��nba5��\+%?����t0�@c�g{�@�T[��lz-k���Y`�����Qʻ�j֐�Ղy�".�v�{H��OZfSdim���DT�&ׇ��HE[���k'�BZ����f�&Іz�ۿU%WNL�����l�F/6_
妒���(҆=�3n�d�й1��V˓o�6�<�UN�uu}Z��IQ�4�0�:F@5䃜���P���y=��kFIr�h��S��Erw���2��N���!��A��d�%�(��٩��яkh���ꦪ��6Ir���S�Q�;8��C���5N���]�W�3+l�tE��o
5�~�q�x��J���p]?bQ?�sf��J������s֍�X�q�}�����8�a6c;��*�T���R���v�����B��հ���+{����<�P\N�5��lT�������燈3�[	��>�=y%�O��L1�x�4��؂�-����[����_�h����9�-���9m�2�Q��w(�m��1%:S��/R�)G�!p�{�ϋyr�j���F�ۨS)��M��mTIP�09�㰋=�o��@k�
�Y��YB�Ŷ��'�g�,�:�p��\�B����ST��0��"��.k�Y�+�ٺ�q�/�>�KBa�!������j�����^�wop�|2�)�e���� 4]{���$
�/�`�Z���"{S� ɕH���&&�^_�*��X�w
ۨ�i4�mwS/c$S�a��c���I��@^]���.L"9j�R��&~C�����s�wyĤ���� Cy֎�_�;�xFڹ��W���#==֔��U��e��)��(�m�%�l1�Qmt�y+D�{�G?��6�\T̪�J��?�+���'ƭؔ�6茟>��d��)N�X �Rp�����Vq^5�:'o�bg*X��R�Jn�M��o�'AAW�`��mߟG����I_�!]����]q}v7���(� ;��0�H��<��+�-_szȵ�i�����O$��=-ʹ��~�4�e����U�)���'��"����&�%<F�� �b��WG :�e,`��5t�_��2)A��q�^�ƠL'ǝ��4�R�C��
!Rewߣ���>]x�(���x��Sj%��^�$Lv�Ѧ<m��m�ԧ� � �&B7l��J������t��+#X�L�_��ʇ��O�ߟM�����ơ�F&�lA2~ٞ���9�$!I1���/ض0�~��@�Ηo78���YuU^s��|_͕��@ݛ��Z6�}�[f����|�hB��n�$�`�D�W0`|@���M�2�~4ϦU�����Ď�
�;Z��Ί㉶yF��A�bi�`������q��\���Q�\��ؙ�u�_�Ɗ���E��������(��h�H��_����QI�O�e�b�|�I]��.t=P��j�
G����Rڂ��m�!7�?�H�d��'��E�>�@��JhC9�R�"�����Q,�A��d]���/���~+��ӪL���N-1��31�$�ފ?�ݻJO�j:o��(3��v��<�t�җH�a�fD��QKج����;Ω��'~Y���G����0��y�������.w�-��v���W�����1�ܡ�O��<��z�,�e��q�y�!6�vcȏGe_ѝ|�w*�Y$�w�S씾�3M�	�Rn�j�&V#L��e�
��ec9��3�ΐ��,t�Z@k@#p5����S�V`I�s��<��*�G�S��G�@�R���y_�W��~7\����e|�|����Lj�6H0�^�iܷ��>з|����B��ZƊ�F�B��YH]ْ>�Q�b�)�I+��5�;6��cY��ޏ��+��wȹĘ]��k�)�[����"���vhOY=��U������i�jI>){u�6E��/&��q:��:\�4�IW�Ԩ-Ñq<p+1�b�~1�RH&�2N�s��XӇ�p�a�$����X���,��d�ٴ�y�	)����������Ǚ��6�u���Loz�����_�m(z��T�l�x3��̻�U^��B��r=�{i��<��;�W�Q��Q|��#���o���e���g�4W��l��E�\h{Xd냣�t.��
rN��(T9��k^�H[aJ@F�6�q�	��p��ܤ	�N��r�S��
B����������J��ww�X����#v��Ҷ�q�P����BjyD�(��w	DL`�����)�,������B>��|�݀���V��J���f�P�a\�
h���kv?誂��F�90�G�����倩��ɘ����-V���k<P����;��4��L;���H�{��PncM_�����܋3u�N�Ϥ#�+���Gˠ��H|��A�0M�������Y�	�a�)Ū���3.��6�Vs���S{@�V@�9"�u��~6]~�_?�N	!�������I��?��m	�ɓ������9`�D�|l�������i��m����Pu���
H���!�K8L]��ǬX5�����r�'.&��|�j�{��˶�v[�'�Ҟp�F��3Ͷ���Ln�0E��8ť>1��/�9�ʈ��O���q㝃Z"i���.�ۨ���h��;*<S@. ��o��¬'��
0¯1���ޒ�[K����!�����:�^����E�VAt<&%�D�b�ˆ����FI��w�]�mp.���b�$�u��_ۧ��âxoT���,��������4+����S�*�6H�3��`��z�ޜ�a�w4���(�_��1 +ݐ�*8��&��� µ���\�]Gq�����O��k��Z0by#�a:�I���>��V6r" �X<\7�4�ؐ���c$�HUs:�<��E��V���l(�Ă{//��#��t.�*<��h��}����[s��c��5�J(���2�$�tĞ�a�� ֘�P�R�1�F�!�{]�#� #���4>�,���
~����}gS�lF�>pϼS�"�w��f
�ᎱLx�N�V0�IZ&��9��#S����k�	��(�Y�c/R�|��dLҫ����Z���ӼL^*4�j��+��-l��V��J_� e��b� �oJ�,�Y�k����,zg�E�&s�u�/�!f���J�CO�����6�=��i>�g�f ���� Jf�$���
��: ��;U����K�ꜣ�0�eޏ�8pډm�];������8���!�=�9�C��> ���l:���̀3���p�f�6��8��<��n����d7Vhu2���������q
�X.J�/ltG�]m�ƙ9 �F���;���7r�[A\F�>c�8�z˰�j�Us�W�`�!*�>38��(�~�������-�qmr8/��Q�|��N��˔�ѿ}5S�e9 o�qDg>�����]V@⽽16`�py���v`|��E�����0q2�[,�1�I�_)��?M[��?d	���@W�R��#�@�!�+=�}�ĝ_Էm�#�.~�@/��P2")���G�ב���u5�Ê>lS3
	����l��B@���h˔	I��Thx�%EH:�����>���ɠ��m�/ ƹ�PzI*������dyj��H̋U:(���O8I�6P�B��FA�Jz���uC�@污SU|����>9
7������}�S'�����_�TP���k�i`=����<f 
~;!���-]�)2���U{6��F!PTc�X�$ɀ�
Z��b9V��ǖ;�m,��w��
�뫸��i��PW�f��p9�{��Cn�K��֪:<�m�Q�qmS���\H"(w��Α���$�CUt�۱�/�9�6^| &��~�9f ��������i`U�,f��~�b6H��棌V;����+�����4�j�Ā!�޸E��4̙Y�Q��7��,�㙕�-<�h�ga��X�x/ۑj��T�mQґ���V!�|S࢛���m]�<�,�9�� ��Q����R�qUbr�qM�5n��hl���(��p�fn�n�S��Ja�����,R��U�_ė~��)S*��i�ǼP8��+�P1�g�V\b�7����C�i�cOb%�$|쪆�|&�s5l���O��k<�b�R���;p�m:�#C��/uKP�����5����M#��ܔٝ� ��ཋ;����^
甝��׌P��,
+m{�Pt�#�p�l��m�1�#:�÷�`��E�o��N+�hU�g�,/�!"����.���Y�r~Nĺt< #��Eb�V�a��h36�?o�H�s�6��qp�uh6�U�!Lś��?o�df}~S�<ϤSOl��'��c�̓0�oͽ�r�wv���X0�Nz�'+޿�f`͗Q&n���44 �=
��*����]mf�:1�FU��cXC��D��vdN���#QP���c�͉;<�Y99���l���sJ�w17L8*X�y;FV���w��h�*���f���H�(������j�nY?�A��q��h_k�]��8K�;}�́� �A�ۑ��_��|uBC�o��b�^1f��� 	�b��������֘`*aJ`['fRW�d�k��d�bF�)���m1��*[8?(v8�,��z˼�=�W�Ća���˼c�x���O��A�D>�uCۜ)�����|l�zw�kT��_�;�9���E� >*߭�T=�H4s��n��V����z˦�b��1	527QHh�.�aL�3�f��IUY��hW��M���`vZ`��h��D3��nG&Țt��� Ӝ[r���vĆ$n��.w>����;����ڣ�0�b���-h5LJqB��IR���⸌C��G5�U�J�7p��ۅ�[rS���_"
P|o+="��L�D/���Uq�]���To���Y-D�`�6)ז����?ra����A���N�D
`�%���x�e��Bh���!_�~~���(�Q3�^������Y��3��,���|Y�f�-����
JwN��It�&J࿁�y�WѦ J!��,��t���/b��UL�̺��r��.��z�*c;'�w����M)ׅF(�f���8��na��P/�#,��?��4%ͩ����Yb��<9�j��r���1�~�"{�n��@��-�cM��H��g��0�!Z6����߻pusj�{����.z��%aY�v�gO��Դj�gУy\%��z�*1u�#p=<\hD4*U��/^�O�9k�2ޔ��z�|�X�|��y��|��|��p���C�^x���(T���2�C�V5�m-q!؂��/;��������)�ƙ:v��yj~.�F#y�Q��@��JRA0 E��a��l�.;6���RK��Kg�	(��a��j�3J����M�����c]}%���0����"_��61a
����%	~��}+0��-�6��c���(�^0.]zE�Q�A��@_�����x�F�����ٚh}�j�	��Vɯ<SW/�y������d g�'����B�|�r��9ul�;^�=�_��U�F�^�N�S]Mۈe#��)Χ��`c鑏�9���i}���y�=��&�?�=y�B��}Y) _���g��b��<��d�P��h�c|���b�z<ê$�ۥ����Kp�uӳ��_��Fh�tЎ��Ԥ�i�ȭ�JOJ��ܫS���f��9�S�rnU�]*ܹ�6/	]U;V	��~�Q�E���_g yx��"a)�^�6��G�-�|�=����N��}��6g�ѽI�%%1��.���A����
�Y����r�7D��2�+��SƇ��;E;r��^L�>A9�,��@�_j�dd�k�@�}��*��,!��E��ɳc��Q��Xս�!�cfY�{�X�&2	@Hrg�0cN�tq��� �ko��w���Tx��/������)\�m@D���>�gŪv�<&�I�[GПB�]Ǚ��X�Hw��c��]V����Rfa��3Q����?�y���%�[C'7oWO��`S�˦=��J}j���W�9��N^�=�}�����y*�Y�>|3�&��P��l���ϰ��� )$-)N�ܐM��Jy��]a��.��r�)C���X���|0���ǛĐ�W���ح�ix��e,5ݛ��YS�X�� �>�?�áӨԷ_��F����ƴ�i�r�BOwܷg��r2�e�hhƨ��<�^Ǜ+Oϝ3_�Q�7󭡽����.��b�@�e������\ b�G�(<[D�"�IM��K�hc�]�$�����'瘰B4�\�e1 m˧�ޒs`4���W�L��=l�S��X5΂�\,�%����}���򄥁h��mg�x���b�C����f�<��a��5��4̷��� /�R��O��3�}���r�8��4��ou�N\S�������&,�+a�+xcJ��f�͔f�VK��7a\
��E����>�K�&C��R~�����G~����zCC1	�f+�"mD�B����kS��*�^� �E�(r�B�b�m�pz�nb�S������pT̐N�^i��G�����dl۶�K���O����h���m̃K �"(���� �Ŭ,�:{��$����X�ǣ�X6�v ��w�ne�����1�fE���kh�b���Ei*�]��Bj���F�P_�o��T����hTg{��I.P����؊Y'gafY���
��s�����J-y�8J�����m���P�Tp��D��z��DZ��Bj�����?G��wǅ�����]9��U
�~#;�`���~��ۖ�ekk�5�u�<�qj�ǧi�߾f��� q^�b��i��'3B!R�?��PVC��C[�t� ���+J�l+�u�G96�>H#
e ��ÇmΆM���|�F�bӵ>�Ʈd{u�q���p/��m��f�r���[g���u�����pE�\�L�5=������'�^��!٬c��rU�6 ��]�����hn�Lݚ��.��F�l�|I�uXN���u�9�7��o��j�깠���ѣ����p`��GZ�ч���R�$ư]ܧ��x-��\�2�4:Lt7Ykx��U�?r0�'�I�sYچ�Z���~rYx����0���L���������9*�d�����ݸ�9�B\�YѸ81e�����eDTA��t�7sX���#a�u�Y����4�?�b����?y�j�*�I�~��e`��G>���v�h����Z72�đ�9~�-մ�LuZ�b���]*���;��e��[�9;�N����H�e �yf��!ŕK�C�o�'-��� -�/�7ͩӫ�:�e�N�������5����]l�H�SCA*BAF..ڔ��ti�������M�@l�g�ĳ-���Z����ίsʣ�n7J��i�TQܘ&�;�c����q�X�In�v5p��= ���iOܰ�ށ\�)g&�A����D� ������K�J�{L���<|�Ӧ�e�ƭZ�g*e� Z�9E�.�<u�������7s.����(�+@��dL �Eʵī=�\
#��l�m��ul��&e�.��	�	�j+�y��{(��C*X5<�t�BxSf a![*����Ad"9Q��c  J��U�E �7qa���J��%h��)���ܖ��b�6Νf���:���%����=������FV�W=��*-���W��l�[�;�@�FX[^"���Gz����ʀ�t�z�w��=z��ND�G��EH᫘(��J5y�-����,���!�܋��87�8#�mg�(�9�K3c���l���w�u`X�)}��#̭��0�6*6��bM����h�瞣�7�7�嚲�<?��t}GAc�'�[{Q@�{���b�k�{��}�[�|�ԥ�0�9��m��(F����7u��YD����Q��>���`��<@� �(��1D�d3B{�0��@��f\�z�0�כ�8���GeKF;2i���Y~�	tS��zk^����߬+K|�G���|����,�P��'Z��b2Mp;xT{�{�o�t�7Ý�`�N�.�:�ռ��G��Y���g�JU�L��!�:~�����W*�)n���'ҟ)��Jj�E��Pa]m.�Ү�]D'pj���P˱���'ơ���ɇ+<W����ޖ�#VI���Lt���$$
x
e�����Ej�A(^�]]q�.��P|��C��ʌ��w���7V�Nkn�I���C���x����T����Z$y�4������/'c��k����N�x��P�23�?v�`İL�
�N�����0 *;��D7ʦ�	+�[q�?�ь��U7��zp.��ļq��t�II���]�sX\��q���p�[�;��2C�N��`a��p���=Z<e����n�8��g�P��JP�)��E}��^7QԳj�m:
I<g����b!Mó���.'Q�J�̢��('�	)|x:�v�?N'�O

��b��������
�v���ŞJ����0�#Kpʱ�qHS���V�dz`-����޶�m�Im�C؂(4��Y�:&�}y�$��R���Jy��N4ZF5�&afg�����&3d��˹�z��?��L���J����A���2�cB���4�>:yͺa}�Г�<ʭ�����vv�,$1��a��j:�M�����T?��vc�]���4d	�^�ޔ�OdvoD�|�˝}=�sLR���_��
ߴ����]oK�c��Q�P6�}�p_=�����n�����)�ݼ�K�W9�t�Q�h�&�t�B�����@�
�Lǫi";�_J��F�H��0�AՁ�|����1,��P���4�Dg���5� P3%����0r�!�[7k���j���S��6/�5}�u@{l������]hE�.,����j����x�
Ep�[�&);��ѕh ��/h�Z[�P��T*1���t�9�/��]�e��0g���W}�����
�/�	S���N��^����F:f�C+MTL������>�9��I�@0g�@;F�����<&�J8ox�Û*kQ��iT�$���������JO H'}]q No�b"9�Q�Q�����?`�J�~y%���a��(W��.n�$(w��#�iyF&A/���Ǟ%��@�Ѱ*{�д�z���#Ͱ����Y�"7/;=�co1�:-�K�6�*ED����A��R����*���!I�b<�©K��w:��;�D�w6�Vd�V��HJ	�slG_��Pv
5�Z���0�Hg��	��3%���lT��!�à�riLP����W#[���Ht���q��Z|�q�$M0���nkXQE�^LB�a0�4���oP��I����B�˃��4(�˗xN��C�z>���|����nr�ɂ̣,7�]<hϙ��,�3�	����m����*�A���y���*}7�Τ�}h9A�X���)���5�:�c��pU����B��Ø,2w�<�=ʻ��
l����@ �䞅���~s:�h��ox��2-�1�,����	�(�*���9�jr��y�c�i~{��d�U����8[�:Da��e���*I`�_����<���8y5�f������1czwm�+���J"(j���H��4-T��aD�3Lr~ws�Ц��.�����d���~Jp�&��Z��[��6,��Obe� ء�
w�?K��>%�bM�	c�c��s��j�;��ϖ%A�hA>c���HM^��#�|��W`4��:k��AL6eϨC/`�)�$�>���ϐ��_� ̥� �N0�$E��/�>)��ic�v6N"L��<��o�V�j�RPƛ���֐^6��	�
S±����b��}:;��H���c���&`k�	��-�jn����1�|��v�Q�K{U�[a�r���Z�������g,��\_T:9A�3��An���I��_�n��=� #��42]m�Fu���e�����ސ�������+#D�e�?����X�GL���54�ٷ3]-��� �'����F��/��}�X+Z�r>�2$mF9G��6C��!m�y�e���2��I����`[�䛒��֘��:0�w���mi~�U��h��!8 ��&R��r����Gn]C�X�M�e^@>+#	x���@�N0�yz�|���h} ����(���� �}b2A��T�|�d.�n3w��/1� 9q��Y��C�{�_�p�[t[<5s��,"f�k�QQģ@-c#�,�8c�|�������d��v�Hm�����7���v�`�R\!P�](��/ϲ�ߨN��' K���w��P)���(�~�D�
n�8��>���i��.����^�X�������B���Y^z�Щ2ۻ��M��Z[�1bL�`.^0�Rk�}�_m?&�3O��]󂰺�W�����N@Q�%{�dT�Э@SG��HM�:����
5��:y#�����#M�@.$��r�}_M���y7xSs8����E��vW�y ��wVDB�閘�X��BRL�6��^��P�XƅÉ\���"\C��^M�}) �3v�Bڏ��\$!�:�xY��x�i!M2(�:���;8*]��,KN 4����2���<R�<�b��8H�;�������~��:��U�t���8��d ������Z$���LӾH�zA�!��_I(����[/����L�<ᜍ���CX��E������>f��nA�}~�� R��d+p�x���	�Jkbq�.�S{�I_n{`1Xx��M�؂��k�~�79zs'�c���fu���;�ΐ��<�c��K�{�ݝ����	#��I_��0�CJ}��ƍ���p\#�9;��}�uk�XUo�ʀ
�jTi��L_��z��k�x�R��1\4�
j�߲�J�v����7���`w����A7p���L���e�
�#�w�t�ɾ�R�Mm�Yu��rZ��_��i��Ja�����vp�'�"`�9�V�+t�8ҩ�aHȀ�*��o���\*Yy1�S��[��'8Nn�)��kt�������x���$�Dl+�X�/�%qjŏ)q$gy��)�M�+XD�둉%���
�v���c�p��^�K���v�(,S�ޯ�V�%N��4!�	.����]�0>=AK���W��~TT��q�n��[�g����4T����Ӯ�	7m`�D��O=��;!s�V��X'��5Ap��KD�Gm���;��N�v�ظ�,0���j�OA͵�>�@�����|��\m��Id���x���יu��jw5h����KY�?&�N�<�ߏ���P�Ԋ�rvŔ]�:���*<Gb���^ �����A�����y
WX�1c���tg�l���垾���\3!� ��K�y:p��"T~��+ۼ=39ͧ������}a�v�6�$=�/ȧ�U^ +{����Q���Cb)������f^�8�z`�5%h5��[T�s:��;S%�i�p~��<E�U�a�Hʈ���5f
��'�
�=�X��'�����;��b�S��~���}��ձ��~��QOuqwl�Z�^�B��:Q�㴵�r��ks��� x�5ZbT�>�iqk�+����l	��;�x�� ���D�=2���u��TҐ�Te�����[}�T�ÓT�wr��"B)�ZP񔀌$"����*�`����)�Y�'򳉄�<��s�s?�o9Y�������˪��QO�e����E�l͸׌�A2�1�Jjo�r]荚�z�җ�
�Y�AQ�����M��N�n���-�̀�H��j�SAn�K�P�	"���<�|7�^�7Y�<g
�
"d����������|���ӫ�AUCS�[���C�{�C5���,w:�ZO໋Fa��#���E�J'Ěs�5�`~({6Ӑ2<6�"Q��u}�U�>�����z�
� \ K�܇���K�l�X<��r峑cmp�.�>��p	����(Y%��Z�"k3�.~J���M��᝾rz��V�ٛt�/N1 ��
-�p'_��,�t�9!���!��K來�@N��X��n����G��@e{�3�b�*��O���}݇�F*,�f��{.&�:|���¨S%�!Od�kjJD�ͥy��NN�,N�Q�b��]��i��C.vQ�2��`b!���!}b��|eq�;}�B�!�O��J��[n����$�C��h��I�J'���i~�������(Í���v�jCw�O!IƊ�ڐUZm@j�q����A�Q����x�XiQb5�|��o E���#I�h��P\ ��e~N����t݆}�t�ģ���_D�ҳ�޾�a��JZаW�Q �!*���:��ܗN�\��&�F��"l&z���`#�I�DUQRm��ـ�Tzq�����7�����c�mÊ��T\��o��$��<iC+�@�lN{X�D!�>D��>���gei�,T޵r�j�$��U
%A�L��?5	&EғPߥ�Kv~Q��c4�KͭX��
Ͽ�EY�M�4ADd���8���$(.f����oD�)��Ơ�:�E�`����L���%�z����j@�AB�0�IC�T��k���)$1���$wN�f�9P����iF��R���F�^Z�H���RwV��ǞTI�wj�O��{��p�p.����6�}|�R	����x��A��tA}�g�Ԯ��A�]�+	��ܗ���r�W�k��Q"A���@�F��	W���o���?)��Ͱ̹1E8]��L�ǧ�a�<x�T��H�B|ԧ�yK��I���E9�&�y�tZ��).����U�_������.ڱB�|?X�(�s��YSju��r&_j�v�����<sXL�:���#�C�!6��=��C��Y��n�K���S��i�v���np�E�����]y�.���-�ic���î��vϗV�,�}4��Fr�;��$���x����^��l��&��L�J���;X(rh������W���]���^�
�P��5��)(�5{��{c��9�q�m��h���W6�[�D�Z�C{�qY],Ƚdއ�^��t�a)�@�0\_Ŗ����-�$��E�,�	����g�������M$p�dG���'��h	�h�J?�'�7{17@���$�vy�>�Wd0n㝁��l�{���D�v�t�:�i��rX)�G���Hb0d�
B\��q/���x�1�G�_گ���27�}���Ư��dl����;A��Yl�.��?�BT��nb�0/w�����9����yԪyJ&,����C}R�sw��K~Pa0�p���r_1q�s5����w���P�%,;bU:��ʒ����Sn_f�鿩:�e�{cJ@W7��ʶ[>��;"��GxֱKQ���F��p�O�DLK�7=BX�ҽ&����s���#�"-~���Y���"�4����G��P�'��̴�+.�7�$��-�b�'0FZ���d@��p&�;�Ο�eų>�͑�����|�E-LJ�������T��i�Ja��]��KxE�*P������+�%�x��&�J?���|��#�o�BES�Ƞ��'����J��������Y�j^�dr��53���L�'G�8�v��חk�m�ⷅ�,ǥo"�nۉ8���d��$>��5%��S>	�{|��i�]�Фj2�yLRѿ
L�A��ړ��ƺF���u�ނ(����\�^���#�?���Cg�8E���p������?�D�!:l� �nr�ΈlAw)�~�P'�Uu�ꩃ�Y6sd���ɒEpp���?L�����Ӓ%���go���(;|��[E[_��3��#(��<��xW Q�*6sBɯ�=����@��/��܎��(,,�^��>�^C�<��� ,U%S�$�k#��#�[�.[!�5�'�����teIt�=����M�����A.#�vc�q�܂5�p��[��	���qˁ���� qq��3��wJ�o�l�}�uE�������Ӕ�,>u`f'���$.mDɆF�:���P ���Mk�%<���؏�ڐ�����kZ.e�(�h�U/7��mY&"��̓�_1�]ۈ�¦Y�7�2$�c��Q,f(^ܟ^��?�>˓;���y�Jn�O���Q�?�cG�k#��	�q&	��\�W�|5�gW��n�g��;��x���$ѣ���~/T�� `�2�$�q["h�t4�ݍcC�w�E�F-Wk/9��M�.���6���h���0���3�Y�*'u�L�$��U�Ҡxh�������{�٘����6�O2t||�	m�vz
�1n`$�ǡ��������,���: a�k���b�w�5p_�\��^�4# AC�p�e��W_8��;K��)�I�!��ӦN�yS����١�����I��i��̔�ӛ�����&��F?�4E����bA���k�E��.�B�|��%��Q��(�`[����B/*a�I[xx�����V� @�OQ'��:�� V�c�����P*� }%��!&Ϊ���{r�Ҙ_W[@�B�t����|��|:ET��&n�x'�6UẍoW�Y�}ق�8�V\F�Q��W3t۠)G�ʎ7mjϹ�mԩ��@aN4�����L�B�D���oSv[?b�O��󄥟����bLV�S�=�bC�_p���f׵�~Z{�Q�ӭ=c�z��ڣ�J��^[�����eJ���R���`��O���UdS�b�i��-#Y+O9�&-�<��ぱ�e#%�s!�:
n=�F����e�[U��;�B�U�t멱��� ��^��������i˟�;'�.!�.�оu��ehaވ���0J]d�c��wv��4�`D�Q�td:��Q�D���T=S^�#�weR�Z��+�>��l�Y��b�VΔ�2��C�Ob���*�#���$�MQ��D�n�?O�����׋J�@%�}WO��~�� r�x�BQz�K$�<�l���u�A���3�����k�h4rW1U���F)*nb�D�ܹ��ЭO/Y�,�g �ZX��T�˨������7Yj�ً�\�}�ީԩ -`���MC g!����!��|�y��5^1_�b��FO���;n&�!�̜���LH%���K���AУ�tE���ȱ���y#+h��Ѷ��<F�ѵ��ЍyR�2����|�q�n�A�����yӿ�F�p��Td�����={A��~��
����k��8N>Թ\.��F'tmH��\��j�1��C�?�pj���ػ�Y(���z�h���aA�Y�>�늀���a�0k�n�2A���(dY���/~t4�S��5��ԍ����a�jҚ�k _8����l�Jz,[��B��gL���J@i���)J0����.�`�!�+�9�L����>�����}#?���nM��%v��MZ�9���v����rJ������{J<���گ����̶��5o��� c���1 5ř&>ōP�Z���*ט���{m r���s�8�߉
�]��7DG������8Ϯ�b!ܟf�1�7�i��r�4E��ad0ՆG�����ecF��2�E�[O �\a��=75X�݈��֟��L�(����GO���� .J\	�凹ͱ�y��#�\N�օ�TB<����s�����eO}�6��-���Fd�E|��U�)�2A~m�؏�(I@4�<7`ޟN���j?�G=xv���`xTO�ۯ�d&)[�	}��aL�>Pf,~v�U�K��;�i���Q��e�@���m6���=<�	K�R*�7���	�Ұ�EJ�LE���.�
i�2�j�U0%1$"�0@�v(0�w
V}z��p/<-�hk�1�19��#��y���w�8��4�{L(���<>y9#CwS,�C��׌�^���<4��h �u��c1!<��S'����b�)�&@�rt�A��>�����Sn��o��Aխ���F�6꺟���"C�3[ �I~5Xg��5���$�d>�@���]��`h3g]1���1�Ri��"���GN�v��Ũ��L
KҪ�U=��>�Jy���ēN/ϞS�����T���
���3�@�_c�%�R9�ҳj)����ߒ�y��W<M�������k��n3��R�ɜ����7%��ϗfq6�<V�k%1o!ϻ�Mè5�CI�2�Q|��Yj���Å�3т�����ξd��l֪~�����p��j$����K���?~�[OF#������� ~�*��b��}��U������%o��b 9�t������(�-�����}3B�Ը:��D��kz�ھ��)*fmֈ9�'�BP�{�&�l�V�
a��u���J8UdGy'�������|d��d/8͈�.��K'��%���U����T���"��N7�W��І���,�g�cx��it���@���$WQJ�L��Ռ��Ɓ]�q�9��QY+}��*��["c��³�٨�ǿt���T��
p�P���ФBգ9�X�S�U�&��>,�s�&DȆI�l����h�TLo��G�`���4 g��0��.�hG��#G���7{�mTu�-V��Bl��X[�O�H?�'�Ջ<�=�P��FzD�p�Q�;N��=��Uo�;��eD@0՜i�MZ�?,�NX����z��8ޢ��ߚ�3:89�A��I6��Ry���Z9�}>P	��c��9 S)��Ќ���>�Y���ht����4��Ȼ?ك�N]�r��[]�Z}>¥G�[禍�	#q��Q���� ���i~�+���e�hx�4&:T���|� �Q+K����I�4Z�,.�<���š�����y�V�٘�H���lz؁��|Y�6i��D�_`��h!:�X���7��'mQ��ђ�{���l������J"�ӝ��I~�Ĝ��]��i7����+>6��%�zuE��2c�����,�`��� �X?��VuA������R�L��K�`��[1�v1�݂`k��t�����PW��q0�݇F��.ǽ���E����*�Z��Hs 5xi`�> ��Z���"��ŽA��"��Mz�i��g_�Uu>D7qۇ�RRYj/��q�ԡB���l���'�C���W�*�_FX�.h�ɥ�&{'�V���D��.���zzƸ�l�8,�S��_ԥhY �%��W �~-Lj;���P�Z�ac$��2�W�٧�N--�(л}d�����,��uב~dT�9�!�Wh��u��<�J�Y��P:�Ņ���E�Xi�{��KS��sh�3� �R�țh�K�@i
A@N�FUAקH��H�?4|� ���%���<L�c'ѤJ�v�[��f�Z(=�^�@Ǖ�=/��yp��	����B�?P�N��>����>�@�U����c|R������yv��>(���u��/���elg�T�v���k���躒��bذ;��7"x�HI��TŌ��b���}yZ�P��Y��Ƈ��n"	`�Q"%���;��ˏ Xkׯt2����D��r���4����C�k�5�U�Մ�N�`��2�r��)%���|ġ�2Қ��>E��[dHNnҵ�~|!]� 7��V�����[�����)(�W�/���?{��r�,�k�z� YC_�Jc�����k_�u�y�ƴ׋�9�#����M�����e`�.pՖ��r����R�,�of��=h��&���-��R(��|]w+���t����<�ߨ�����ttk!ŗ�����AҰ��c�7�:w������!�{1[f�T Q�M@��{���PJ�|2#,��-*/˓3�
�y�vH҂d�Y���]Jo��_&x�U�����#,��٦_�H3����x7g��ro@b;l����k�Z��x<v�c�o����pk?G����껨������m@.����j>7��ڵ��$�M�ZD���&*b H���ml�ym��1ȅ�0
�p�ӡMy�f�z���bnS����@,�e��
u�:���ӡj��Ci��wVR+�WMckC�����\��BlH�@[�¬s���x�~��r�t�t�����a�Q�zk�C@��H�J��#���.��׌QUIU�������l��b��o�Ttr`s��mF>(N�&��/�V䏗���7�O�����%���7µP�6��S�k��_�)����.MQZ�<��'Rf_��ቁXk�ġ:���Q�p��\;���m��Zb�¬�,�|[ť���r�Yw	�Ca������@�8�!�ZF�+/M̏�nYR�>u����������h��E̬��:��t��'e7��^'��my��A((�uEz�	_F�)�a� $CA�ӷ@�$ZE�Q����O&������-��<���sK��p��,&}� ��į�Е����z�(�R>��_�F��9rg� tm\h�}b�^T�8 � �$w��
sJ��㼣G^N���R���y`�tE�����(	S����8�d�0&����Ո���{����p䮗�QT��bҮ��i�ڭ�i�����{��u(p�2�3�j���7En�ӧ�F&'��o���)���c�����?Ht�����A�D������tv_o�h�
�����o�
8�m��r�EV5�'�$������m�K2��ֳ�4�ktI"�������ė�0�菦��k�sI iu�)��Mfn)̒7�E��?�<�MK���>ӵ�6��Q����'�O7ů���\�P�$Y�Y�~����b]"�����Y��x��S4c����g����~���Nj�p��P��Qʌ@�<��ض�Lvk�z���m)�G$�P�ʋ\~��o��d����15b�0�����:�:�Stvh	Wsbt!�O�\`�1�7����'��E7R��4(��	���3Q���b�l�]�fs������W�:��,�Y��SEe�� �r�zb@$�x�"n5��.E�H�^p{���je�@@��~.�<���L�ޭ`-1�ɀ���P	n�ߐN�3X�堡��w�ҤO���[��f	/�ߢL��Bن��i�ݷҗ�S,�a"��r��A!,M� ��!�.#�?���d�Y� j��w�k-�5����z	v�D���\��:.##w��F�p�n���&�WHl�C�=jm�E���Z��#�{�q�-�INY�ݍ	N=@��{�ޥ�4Q=��2I�Juk_r. �5�Mc5^m��� �RG#(eY5�k�6�!�챧=@��j7֝�����|�������$K�Sc=5u����LeiO����6\�̖�s^*�%����M����5�ǭ�� 7h�h^���Yhn:G�2�N%u2t��C��lY�Ρ��@�#� D�c��7��f����ǀ�pR����i/?T#46��ջ������ؒ5B� �x|rz�g�P�Հ5n�U�S<�����v�J��Q�/�l���W��v�8,��<�������e��'ܜ�ċ^P� Lw�_��k�%F((��&���
��E��_�$Zбw��� �-��o�=��� ����oqm�}A7���ZK���yq�5N,>vn+�$w؎���Cw�2�5�!�����ҵ�//�ڽe��jù	M���^VKd\�l��L�_�i�;�/=��VOd����ǧ��2}@S��S۳�~����i��z�E���ܩ�GԞ���gR��Ň�>�{��z G�Ej}�>��`4{{�.��9���pc�Py��E��7e���Vlٸ��O�mɄ�o<�}�ߋ(�]��U�����a4N\!���v例�z�3�;��w6p6��8�"�M���5�(�W���5x����$�*~�]Y-�]���2w3��|$Vò ǩ�K͙T�Yⅸ�!�r�+p��EJHg��0z�oe�y�m�ǁ��&j�ĺf!��f�I�>��`0�{g���؜�'��aQ��p�[ק>��B0k������H���r�%�VI��G>�QJu�����o�`mD�:^�~�0I���&�&hK|n(x�ap�,���L���3e#h֥��4b8 �hԔN2O
�@YܟLQ\:E.;��:Ӛ�q^�x[�]j��b _�����+�ݫT�����Z���+b^c�� ��YǓ\���Gq�֥<��R�_G��_�ܧ�Y����|�����V��I���ffL�F����j]���1�#�2it�TY�\����{�>̂�V��>מVg$��VQ��w���%��ĵJ�E����PZe��e<�,6���|s��Eh��$ԍ���-ϺpV�Me�B8�W���]k��k2sc"�8���F7��u2O(��Ü�m~�H�s5 �-�]��X>[���CN����r�������U�'Kr+��r����E�GbB_��V��v��j��� ���2jd1���(դC�c��#��T�^XT��+�p�(.�в\�2�=�K���5{��P�T�r��N
X��S�u ��0EI0��+(���>TB�X�|@�C���P�5׷)x3t���T���������\�lA2�˚k,l
�=�u �.�P��*nl߽��8��_&1&��@���*5�Jؙ��p�ધ�>�?��q��"�1/��Vj���{����<��:Y;������XFI"&�3�00�\
��	�"u�`�b=��\#��l ]��)/(k#\Tn��j ���MT�W�x�	�;�xA�����{���'qz�2�Q'4�^�|�L1��"Z��!���NB��! �V�dʆ��B�>�f�����EY���z�ث�����$���K����ݿ��O��A��Ɯ?���<��{ё�� �+��Ѩ�����Г�UgI̙�	��J> �/����۬U��*
�x̥V�?��h����/L	H��Cj��[��RG/ z��v�����)Ɇ�����R���+�8�b��`E�#N��@O_�1�}��Zl��C7B
v�Ý�����"�n�TxtU]݂St�s$��2p����N�B�٤j?���=Ĵ��8��nH���} $����t�,�l" ��%�=��ތ3���턗�a�~���{�C�Z��e�|��8Q���9�����^JL�$�6�W���p���c�S��Ê�l+C�ƫ������rX�Ax�_�Oҫ�R#;�!�!������LK�fi���ٳ���}��_"2��cSyj �L�~lR�{Y^�V����A���T�%~n.vϞ�$2�����>�F!v��]3~ƞfr��?Q���_n�+��b���Yآr�-��_�3�F:������t2};��G<��?�q�H���zM�x �K�Ћ��5�ގ�rNl�_,5�2�_YvA׵�s��,�!��s�����>�ji�϶ەM��'4i�ah�j$���r4��H����C������-|����(?��m�T���)���6�W=U��J�G�ޮ�=�q�tL�j�y(�b��F���%�vk�ܲC�����O9R"~`�KËH�n`(�с{��M#�� \P؛2�d�B�
�F�1W�rD���4�A�7��� �(�$��.U��m#��y�t�8�`�d>�3�}����y�@�.�X}�B������&Y�L]_�/�|�0��|�dp]�!.�ɡ�Z��KGj%��XC�	TM�s��'}��c|�`y���`O�V�=�g�#|5aħ��MPi3+�_(@7²I�?S��A�-�����&7[�*_�K�Rg_��g�Y�ӕMk��8g��e��8̿|5B-YO�r�Vm��rL�D����k�d�h�z��
yT��w��B4i�?����O�2O���S!��Q��K�4�x�o�P<(EoE����H�/j��j}��q�[C�C�N�^ d:�֡Q@���9�^T�̞h��u�|>�p���1L�MT�hI��Z��,���'=/����2�t��*�W}J@'��s��4��A�I��[�i�,ѵ�6p����c�A�X]�;��?|�r�C�1�/����^׾��������<f3n�(�i�h��N��������/�����߅,�(�Z�{>��%��ˀ�$�-���D��d�O/2�*(Ko��U6BK�Ĳ=h���7��d.�QH�̟9,��TS���s��-�R�i�⽯�������$��Ȁ��U/��� A9b���2�**y�Ɇ����b(�9���l��2Ю��JA/:����I�X��N���w�\@���5��#N����PyUZ;/�켯��$�%ȶJ�H[�����Î������L��vi����W�<�)��*;4�0c�=�R��Iȉ�zY4���-���F0��##��i�V��W�@տ��h�Gf�mxu����W�����4���aUP{��Z��/������xkZ���8v�IP�*_/xѥ��v6\�a`�E?!}��1p���M��h�ɫ!�{eS)�y���M5�#�,�8%+��	�u��=���D��jΆL]�P��3�f���	ml�I����ӳ�
�g>2/����"(���}�6�{M� یZh�����+,�l�T��f���+�0��p��Ue�oV�!+D���)A��2��@�Ћ��"	Q�k�̎��	��N"�&F��V���T��v���{|������v���2�9%���u�C:��;�b�꿩R��R�{돆��{)��B�Bf���c�_L+�7��~aͺ���q%�X��ϑ;��=`�)��B���J�H@��Ë�k�0�Y�����</ޓ%jU��o�b=5m�y¦��}V�kt�w�R�r�_�h���W�
 ��Ikl�s��ҁ�-�ˊ\��?П���+1���מ�C�'�w�q|���o�X���y�UV��8#\g�Z�`�˺K�W�x,Z��� �:�Z����cC��m
+�BJt0�d��	�=�_V<�m1d󇬇��?Q`�5��(G����JɬFM�9�Àx�+�՚:��8*@�|���Т�Zqz<R�F�c�{�t� V��~�2�.\�C�$=Ї�X�(�ŧ}�3M�n�O��߯�*f[mZ^����q:�l&׽7�=��ֳKGs2���q�1:"���i{:���xc_�3�ҐK�ӳSxy>�d2�pCXx']�aے�Nw]�-R��c�c~����t�}D���;���OH{�b�<0�C#}�]��7
�n�+��R�Fv����4K���Έ�4�}���h��ͭ���W���L�A��Sޒ�f
WG鈔(B���g2U��2���,f�GJsTK6:���!2�7���yy7����l��e%9�)K��%گ� ��0{�lL���Lo�ƾ+`���c-�Մ��X>��D&��fR�aΉ['�\�Cj�zV���-\]�2~�r������<Ё��y�8L|��|"�k��%첞�3�O9�21D�&���Y:>X~S�·��W��'x�d�n������YTz�g�C���W�o�E����hȣP�9W0���:��N��%��+�*t�q�M��?�����%,�#9;M���:kΪ�<^U��N����B� g�,�����"��>��M�����,>n鞿!�@�?P�SQ���F[�x"��j�x�n+�{�e��DH�d����C��͐���/:�z����J	�0G�w�]4�j�1�m��B�3n�t����7�a�����LKNe|}* �u�>�b�Y��X������e�p��UA��HV���p6w�j�/�*ʗ.)�[V^>S>�t�����m���^tD	M"�X=��C�+�h	gW;�^�]��El�Q\�r{!��v)���qc"��ڴ�Ͼ��^we�G��`i��ՄQ7�7����(S,����Ð	i �e�)W$�e���\����P�T��X��X�M/'��d���x�y�ǚI�� ���d��SVH��nD��ǳ�O�:��u̷涸�����w�?ʙ��*�e�i\tW8�8��+��#��G%�Y�`��X��.k�{��m��*ü=.%O�?��UH��ޕ���
�H��Zm#�d��6k��V;0v�����j�>��=������^�M�o��vO��-<`��+���8�"����P��)aT%�.����ϛ�î�Ä�dE����u�7OF<�_�y�3�`ŚG�j.��z��`��t�N����$��VU�i����$[�ٿ�I��� ��:�dO�J�&��X�U�0���!UL_9n�A����f� �&�q���*Q�%i��(��Z�Mp��aZ�m0&�6b��2��g�z�J����b-����)tq�o�p��?�ݥD�N���gE|k����H�)O��hq� IE)s�d����B����_�v��$Z�g�?� 0�K���V�3�RŴ��a�K6���L�B>
sov�3�[����܌aoYh���b��S��*"57؊�@���5�~&�gS�.���j��MJ���i�$�x~+	��i��\��r��iB)`.����u&��WT��7���19b���w��j��HQs0�Z�O%�ä�g���:�����{�]Z����(��1A1Huo����9��Qa&3^��;�Œ��#�r�D�aC[��m"����G��#Lȶ q��V����,el?�7���ѐ�\ʩ|�Sx��gk+I���:�pF-��	Qc�� �'U.�{QG�� `�S]l��:8L+h�R���J���<�QC4lo'��+�;�v��!�
�p��/I������u8���|q�W�D';�>$
�(#�b�2)�Ш�pV�x����|��m�P�t�q�p�/�H��u)��Th0�����2p�'��*$��%�ِ/�Hs:�-�6�-ښ��ם�%f{/z���D���Mŕ\�&�P�
;��@׃�j��$�F�!gd�SF���Ehk��շ�yB"����Q5�H��Y��kB���M������y�o��"ezOJ�F�m~�����s&9����C�q���ؠ,w��wh?d��agV�����51��&ZOa���GcM L+Օӡ��2��׮-yOnY�� �PV��C������
Ԗ~���f���Q�[��đE6���uۤ�Ю���@����x��s���N�T&Vn��}����������~[��}���d;BU;Yo���e�	a�<�y~��3S�t��3~��§�M���9�;fo��|8ƻ����H|f^*+ۻ�&ߦ�-L����J��������jO���=27��좛ل��ۣ� "r'���������I��L��0\i1���Y!��:UȈ�tPsg@�jcF�=0KˠgD1Ȳ, �I��[.;J�V���H<�;�N�^z�8=���m�kq�q;� ��!�&}�A���TpZ��'���#�Ԏnf����$֡��/:�"�2����>������`����*�㗁�	2���F���I�__��oas��a�E�a�It�[�9�4�	QX�ccB�4�&��Ж/��d@�XH�	D]��`F��79Z����F�c��&�芢�0��9^�ڻ���<��\]�{���� ~�܄wI��W^@I�Nu��v ��9��:Ɉ�qZa8�U�i[Z��J���^�4ލ�V��`�f�����PO[��ڄ)y8�#�#�s��ɢV�����E�W�ڰ����G�
�z(�/�䏐 ��3��H)�^s	a���:'4XRnoS�gK�Ozհ�c-=�yCɉui�F�,
=�V^M&�ni�(��2|;'w����f��*~a+&�$=��@��wO����p�	�^M�Pє���wv4��W���Mڕ��A��"L�ʼHz����CQ��.@���S���_8rE�	�^0e��A�K��o!��ghf����t.����q��-���C��GE����X�h�%j�l�2�c��$ƴ�E|��� ����Z��ui	������t���k,)/+�&�v.��$��9�sU����&iN3�Q���5����OS�������Aa��j�Ґ�byB\[p)�߃QҹZ�0f�4���B���j��֭���3W�u�?6��y-[���;}�6�6���Hٞ}z�3z�-`7x�J辡�Z"M��d���L/Ƿ�j=%�-F1��Rf�{j*ȧ�>�˟��T�|�B=t@ޘ8Nz�>Y�v���������emF\�)>��œ�$�
='��<]rK���Ŏ��5H��6�Ė�y�'P%?w�,[���u���ņ���'��3G/������2o�Cӵ�R=7C$�F.���*!}���7H��-(�H�H��� �=���l�{11���=���(ŋ�b���`���1b�Xz��5f +��������~��ǽ!�Q<8,Mt #$��X�ݚ�1�~�2���+�̯�s�ш{P��]�&{%6D��m|O��]fb	1VP��y��>��BE׼�� ��*������OIX�W�\��s��EF`�An$��2���a�A�I��r�o6N8�^����bf�Ջ~�T�פ-�a*tw�K�E���f����@]��[���"j]��g�J����@�Q��,��(�� !�ƣ5)i �Pol��Ŧ�Z0tve�v+{E����fv"�r4s����l_�j�����2+��y���o�z�?^筲�_����,��o��k!T(��Wcd�����V�h�$��e�L��� ��o}�ܸ%�͠�xdW#�(�Ů��}u���<L���g�$3�oGE�U�
�`VF�W��v���Fa��*��|�����~g�����i�zƹ��Ĳ�i�Fw��.a:��#��!Q��S��V�o�p�lW&ɚO��#�k�*vjQ)��R�sPs����8�9:�R�N��)�&Z骱F�+���!�����|V�D�"�O,�t����uq-���y ��]��T�@�D�w^�Bp`!
��i������>����nqI+&4��=Fq���\�D݈W��P���r��X�Y=#V�<cP��_��4�H|�v}��6���z#�T�w"�Ϗ���u��?���$?���\��^MK.����!��A���p���ᵏ"	`�5�K�{�(˫�S�d�1t��e�i�sy�pȆ�:h��
�Mӡ��U,�m�8J$Ysn��ߙ��["��R�8���v%��-��w��'�R�JN&|�2�b��-��-��f����ܜ|�>�/�ƒ��Zo �L�R=�A���N��ND&٫i�2^,�3�kj��~� ���d�w�t_��9Q�9DmP���4�hC��߰�>���(�Ȕ����F>���CѤQC�,�<�`8z����-eY�|�#��hR騅���� ˤ(3��K!�:zY�1��%�m�<_�x ��{�E��b�?�0?Kw�ښ�+�`�\��ә���T���-�Ο�,ʲ��#U͸�|w@"w�+S��p��IM�bK��G�Z��\�h0�0�8�:�)�ȪQ]�3G+_�=�d�[m�0�W�N�j0J�v;�~�I��C�8�zTT�P�������
f;��P'���5�
\��(�V��1cG�����T��7���+9���{!il$�U��i��G=��� ��� �n�y���������AT<�"�̯WL��8�>%�H����b�F�i�B[�c��Ktmy���*�$:���Pa�9I������t2�݉@����8-��DO���zl>yI���Ow����͠e3V����e�ѡ��g+�Эa~������O�	#֞�^rغ�z���o�vӬ����ʤ����kF��.�r�-��.�b"�y�� �(���ӑ�yXH:-ۓ��c��~�����Hz���������PG+�c�_Z歈F�a����_N�����fqEM��D��͚KC<F_�|�8�({U36���7�lX)N閊6�p�>���p���%-e;�L����&^S��k�b�g���Rr�b�~�`�Χ�PX6��0ɜ������kg��D>�˚~�[���\<2鍅\�K��Z�  H%�t�N�&`*,>��9t#�:��
L��"ȕ�~n���\,���	�ʹ._���͹��4�֊ZFٮ����+��{��kv�d~񧚌d���TϗY�(3�s��D"��VϾ���p���j�N+@x�H�Z��1`\�^�L�7�R�+W�؇���nI����S��>�����v�#0\g�o���C��h�=�z'�.���p~�/�NIx'�� ���ש�s�9�HS���w1���P�RfX�$��Z����,���>�7_-��O=;ԸΥ�Y)���_u��$�ѣb/7]�~��[H��wԓ�T(���4X�"��AH��Y�QQ��`vl�2#0L,��Q,R^��8��G\�H޹1h2�
�<��xm�Iա�ǌ7���$���"����u�0��+.z����ͥ�hbT� �.���� ٯ��E���qP�Wy�,�&HF�K�Xڎ�0�"��;��K�-yk�ٲ��M.?��-���!+�w1\��G dь�l�@Z_u� �4V��4�r�R�G���cW9���{	���q��(-7�؈���wd$�:���B�0�[���l�G�	�oS�dn���սc�8K�t�@@|�WX�xaum^��|y��3�x ��&�`��p�R��^惶�4u#XN��x��)����@b���@��۹���y��+���`Dw%=
��+T���By��s7�2?��/��1���u�7.�C�^��`��8�~W��:R|?o������+m�e�9j�]19��*d�Y<c�i�&їk�S�R�SJ(���;� ��X���ؽng��&��`iw�����T �)s��ﰾ����K�'
��6*}�r��@~�������3I^x���yd��}#0)"�.�YP	����}MT��Q�l@	���	#��}	����t�f�⤈�/P�Z�hKR[R�H�M�u����Ӄ�
���U��[^w�4-G��Pt���E��S�I�ˮD�z]Nc0�9� K���o>l��o�"�9��5�̋+��1-���z�wQh��8|͖ i�$;X5�D�޵�G�F��M���r�fs5����R�@9���y�9�*�
�\f�t���O����J��٣��@��G���,���5Pmdm�ȶbX�M�7����7�=����CG�#+�d!�Y=@��ʾ��X�"	Av9�2r��"I��?��o�:a+�Jqی�{�1�o��%��S���-����F����ݛ/�	��і%��$�2��8�І2�R̡�1���r�M/*�9��2C��\�_N3���~���7 �O8�%w�X�V+-;�Z�cT��$�Q�|y�S���d}r���T}4!,����8>U(t�eh�F�YnT�B�RQO�@c߸ e��Øz^}N�M��N �v%$��Kkf	 ��_!�S���FV*"X$Q6f����#�.������ ��fn�E)U����{���U��ޮ��d�_��]@��E�����&��C�İ�����G�����)����@�9�����w]<y�~�!�e�����BX���cNz��ׯgk��[��������xQ�l(�}�Noi��J����<��M�k�{�2�u�*�U�7{�����[v�j�}���nuA�vl�����(�_�S�&o�zP�m����]�&�S�_�m������i�-��*d�#�ܹ�т ��bGcȵs�,�d��:YJT)i����p�򜆖 i~�;5X��G1��U�P�'4���ȴm�]����K{�Q5���bR�������q���[���@sq��-�u�$z��I3��H��ǈ����+~F��¦=Z�$�������>��f�-���� �Y���^M�j`eb����Y��)NZ��Z�n�m�P��Rr�J�����i0��ⅳ��Q� x�IB�h����w�rH�X�S9��d�����iǤ��:0<���)m��"M�Ä��I�m� �oE��'�����[�"��EX,O���JQ�7K�!�.Y��)�鷹�֜��Sޮ��Q����)z��_��)�1gY��?�}�/�]��ެʻ���GKKe-֡eG��ŁKr��2� �V�k�*��m��O�%��������1���cP��gnz���3Wz`'w��;�|�N�)0������MX�F�'l�=!1��7���Y�e���`�+$��83U kŎj���N$�M��H��U�8[�Z���.ʀ�^Aa�iZ������x�� tWŕ(QQC&���V�kHB�����*�=�����d��F����-���SL�T��{�����Q۷f}�w3�j�z���8�����DJ[^�4s%� MA�7�X��>�	H0t���#Q ���sv��k�\0�f�J��~<�i*��r�3���!��@���W����+��FajAd�oy�7�!�AU�9_}�1��G	�BeNL2@�O��8����Z������O�u�J��%�qQVC�ql� �wc���@HzQ0�~uqZ<Ne����A��3�-EԀ\���	�;����#��6�/�sB��Ҿy�'WC�� `���RŻ �f�̷�C��j���;[Z���~a�4��qd�r�Bu�g��֯⴨�O��T�);+�|�X�R���Dy�#ͱ��x`{��������`I*�eͣ!�}�z<��U�4��v�����eJN��&P�-��^���ݦ̽�����=_��X���~��v�l 
֌o��m���A�-�y���� ⢛�$�5Vh�"���,�1�ӑA�0�|���19���r���(�z0�}�+�{����m��?����mL��!�/��i�t��ѡpB[&`���+Rd嶪�	����0g27	�p7�����(R����q釔+<���m�N���ެl0d{&��B7ǙG�/]i�l����(;�8 T������7~�~NXP��
0����H">�N
��Yϐ)�I�r]By��X�%}IJ��F��S����f/�h�Th�a�Q\�����Ͼd�J��)���CX�x���dAV��=W�n:�g�?z_k�� �ބg5̹HÕ[��K�"3Ȉ��j-yω�J6�Ĝ�\��y
��%(���R�G������u{'5n-q� �7������87� ��E �)�d����Y�Fh�9&S��>�Z������d��A�B5�ȳ��rvLkŴFj�",(x�^ϸ��kmI�c*��[��Y>�/��y�@�Z��w��lG��B�>j5ڈ��fA�y�g�o w��#T&��;�:��U|�o[ԛ?�ޏ�V>��:��r-�Uu 3Ǉ��?|8���ƒ�7�{A��� ��B&�ߩ~��P������`$���X�)?���{I��jک�!�mﳗ6y��7���n<R��w��6�R���)� ���Ј#$us��
�7`{�x�Es���=���;����JʮJpW�l7�
��+�!�*�>~�]2 ��z!�o��7�>J�	�����ˆ�ʚ�C»���>% �5t��-��C;v�n�Vd������~3��~��/�  �q����Y=��I�ۆ8�|+^u!��h>R����So
Z��%���;���o���K�|�6��O�*ȴ;0S,%k�>���q��L���s!�˘Nc�&oy���_��܆�[�`ǔ�a��3�c]��,��I���!���T�NM�0�;�q��f>:���6q���u�O�F��&��i/�8�̺�oM���(�Ct�S���3le���6|��N�m�u��hB+�4G�Sy�q_,msЫle�[�����:�2�V(�6����j�T�4�ٓD�H�j��+>F	+�7jt���Xb�6�^&
�Z��~�hD1IQ��퇗����G�X��"������ -dH�DfX.V�����H�%�O��3Dg�����[�	���γdI���B�Tꇭ��]�1�Qȅ�ă��o+�%/5�(NLOܚ%�����H0��z�x����䕆����B�9�|<�ݳC��X�$w�	N��U'P�J���>����P����@ūX;� 憥"?�l琖^%�1����Q�)���v�,�g�ږ�$;��m�ga�fl����j0uf'D�8����D�Q5h�1k(hLu,��,�4�E�6�|�I�"�f�S[���t�ib��e�G�	�Q��,kl�1�Y9�=	FyO*�@��A4[��LS���T��/H�[���/!s��8
1$�Ӥ����6P^���vG�p%��QX��t��rs�����5�#`]3U�w�\8��yz<��Xز�|*��t���x�M�%�'�b�y�5��Ȏu 3kd�ndq��ϻ�+�����X�����|�� Û@���סt2$;`l%���`��~�Q8'Z��My���r�����bxK��sܘ<Q\m]�0�d�X*�?I (��݃�,�uY����RY�o1j�zq$����4)/��Iߠ(G>���NuMX�w�r@p?J�_@�8!n�ºr�����Y�UN@��B��N�r��&}t����J�.y,���{)��a[���g�E�dpF�D��G�7s��!n��އƬ�̶W[��D�R����^bV�s���Dgkf�����"�Y�����"Swn�Mrn<4F[k�Q���ӑt3w���CG�53��B���C�������H4�?U��~��(-�;n�q�	{�nut /�<���Ҭ�)�PW-QD���Ҟ>�.,FF�T����#\:�s����U�X�$�+��1�"^����� �����$���L�|Gk���<W4��@���7!_�T�b�\N�	�X�^_	Yw������~W�'�L�$�od�<C�s1(h7�4?��V:G7��,N��-Wk��k��^)R�����,�W�i���P<LM|b����u�xbVt"H�Z,TL+EG��U�J٢�"����k!	`��+q2���Q��j�d&�;D�p,0�?�MI�`�`
Cc�ݰ�<ɍ �}P:�(+�t(�-�{��V�YY�+��Y���ۄW���MJ��Q��K���_�O%VT�nCZyc�>�o�>6�Әа�-w>x6��X9�2qQeM��ݐ��m��`�^o�)	��X�>��x8��GaS�4F���\���놌�Uө�z���9A�/�ײI8ph�NQ:2T^A΄5*AwH���3~�_�X��H-'�T�o��k�0�ް���y.9�B-t5T�:q%Mum�:[�3|���^��)��㐋��1��wR"c=�:��z��hs-�O�
���[>�e{,z��Th�ZS�Kc��]��/N�ʞ�� e��ˉ����ۦJ���1ɒ�v��D�K#w,Y@�İ�Ǖ�܏6L�嬨m}�2��q��(@�^K��f�,��$ټ����/	����#�xS�~��$V~����*f�<��Mo�ژ��3�5�ܸӔmh�~Y!t�3�����zDCc�W����t@�*w����uP#��]_�	�W�?��%L�R���މϓ��fW+�EU�1 u�a��S=�c?��BC�4������,�(<���L�B3��?y���s"�U�֏T�+�o��מ�ya]����dբa�u�P�#���Z��k��ו���D�ܧ��Ө��:���h6��p.�8��ap�.�$j,�K����k%-Õ�$���{ԂD�������<;���0%��[&D��MĹ�\c�S7��<9S@��A�l�$Y�}ʋ�wVH�Լ�Z�3����F�I+��N��r���Q��2~�2�R�6<z��Q�a����T1�V�R�4uF���y�����=O�������}��,9(�;/v�K֕������6 �Y�S�[�9�/����Nr�0E����S�ǹ��!�9O��I$�8���sU�m���11*�H���|�X��ck,B�Ӂ<��D$���DrksJq���ŀ�kD1������������goѢ���咬�$f0Ml�S�I�4�H�L�ID^�yA��.�m���"���Q�I��Xf?JޤJ �Ⱥ5 ���\|<�ݕ�������s�d�8�m�zg��fY��V��d�ȑ��`ui?C�*D�ӎ��O'_"�^�Ҿ%�y�\�E����S�h���Q�-�) i:�Hk��y����s�At9g����1�Vd�ϔ��^?��T�����Bw��ל�B��;X"3@�|R��>��1�o�j�	<fP!pdB"�|��<q_gG�M���b���oy@T���D�rj pФ���j�_���[ۨH83�i�2���%w���r3gt>�@yNU�\��Y�[X>X"���VVu��]p�1I�@�x�}��w���ZR��@�n���,{��f�Z���Y�ӱFD��7�_�{��p��e�`����(�"�-���H�H>U�szͲ�q�0L����0u��&�����T����b	԰�c��?��1��&.�[�A�B���"�WqB���u���[bƿ���
lke���`�R��H�b;{"���o\�P6�\�b��j.��S�:��)���7P�����MUZ9���&�a�����;$}�omy�?��__o�푵��z*[����_�,Ț�f�`FF��XS O,�DP�LԻ���SYn^��?�O$��O���G7��!�烖",�^�K�g�g���\傅���R�p�kV�
�ϼ�,,�K�<m���?ߛJ��O��c�^@X�H�Vq��|B���5������C
����f�[��3�.������q0 o���X��?��d5��2E������d؃�s_9�R3�ɜpVQ�|p��#��C�'S ��7��TJ�4GP���1��Fe���		.�	������z�:_��D�.R�DEL\�׮�b��[P��X_شT�K����2�n�/�V�Z6�y��.#U�Ӫ���%,.+E�V��x;��w�JQfI-A6DC�]ʐ,��x,#���c�{�����2�Ή��1��3[�GɮPM�a��]]�1�B�� ����� D�n+�3�@Oċ+=�{�C͋�t���K^s[s#NʕYYy�>�iM��;��I*��*�vߙ9�p
�v��0���f�֍�5�s�OF~�=�+�RUD��MR�^�U��������Xl5~�;oc	x�E#|$�|�1�ǙE{<K�����/"T��C�	��҆S)94ÏB)�:�Z]s�J���xWba����wM��r���Bo핯>!�\������)�C��3{x
0˥�/��ĚD�6)�eU�A*|���w�&4ŉ��Q_jh���g�����_$�������o��g�r��M=|Wu�t��/cLN�Z�I����$� �Խ�ua��˔���{�JW��"4�3�B�8Ш�S�]��L�9�{����}�Ү�{̼�r�+���^@�L�2j+SXGݧ���鴃S���|��K��=M�'�k�.� �SM^�r���D�q�8!6��QyNj"c�ø҄IE
��V�l7�G�à�[�����'����(��LG��<Z�d�رa<��2��
��H�,Z��?Bg�dy��2�N��t�&��&�5���4�k'�6�5�e{��H�M�;T㙇LHu��̕�(���8�	��
����ʽlH�xL��"�t��!A^�x�~��{�d�8���D*C�Y�$.	m�9�(g7�oP���v5e��oQ��w!�Έ�q��9��	2�c���jԄ���fX���W$#��	i.
�v����I��B$/O덎��9��~�^��V2�J0lP�*]۩�q����e>��v��u&y�&6kAT�_h��G���AY�E�	13*o]lK�]�����H:q��`�qኁ�#�7� �J�ڠ��;k�?@ܬ��w��W|9�|F]7a&vz�V����&��!	!��Rl�&8�W�-gS�ĹO���V��v��+:������)^�։&l^`�D�wWeZ=��G���]�46��K�eo����®��	+����Ǣu�C��Ԁ7�Դ�TR���T79�ݕ�;��5�O\+HcE� �*A�+�=.���Z��ŷ��JFz� ��iD����
5G2�Xy����k�F�eoiԳ�%�*�~�.�h�\�[�[�@F���x��#�y힌��.�^\�Ӓ�K�O�x,��Y����h��mPQ+�X���1�.b�B
�b�;��_̅3G4�V��Ø�A��{��.�F��*����6! �U��Ϥ�t݇�|1��I��_���yiB��� �yDy����Ì��Xt5^pB�������z��m��u���g���W7�ǖ�T���\fs��f�F7�����,�ͥJ��#�^$A��v-9���S  ڍ�"�g�0�eԤ;^̺�Zړ�dF6�=ldK�?�d��@����{���ǯy6�:��a)�p=-�_�_�[Ψ2�V��Ci<���Y����Tfy�ӗ���	ʑ]�f��K��@�LZ�ܖ�DAUUr2��6��_�/�_ʟns8���!��YY�x
k0��_��*�G6��Yj~&}�a�G�)%
z)^)�\'�)��F��ضj���<5��-�LV���=J\N����!4�v�L�坯�&^�~�	�h��.�j��΢ڼҚ6X����6ɂ���5���Z��|1����v,m��Tif����o��<��������U��3T�Me�[��M���y�����~D]�wG�y�m=�@�3��+�90�� 6�<�WG�\176~r�a]{V�\4���۵��UZ#�g��b����̔;^>;[%,��|E
�J��g�x�1��R�z��|\ʵL��uL��2R��={+U}���8&�) Rk�C�������r�w�SĀ�3�"�Y۠"[�=�T�C�
�:���ì����ٴjt<v�:oO�k�A�v��/����D����6"�=o�M$+����x=T	��^�O��%a�a%E� �ÏyI*�|7��w��Հ��}%�q��Xy�Q��@a����b��4��� �_�w\��o��OɅ�Ũ5�aq1�r�T]���`_��@ S���Z����7$u�#tr|g��%�Q�����m��OI�y �꽷~Ö�`
$#b 9������(L5"@|�{��1@�"��mN�N��F%w�y}��R�����ۑ<��qJ�y9@��j,�4���,�y"�1���ߎ��k���{��:��W�&��	Z�<q�
�<�_��tuyfng�k�
�|2)aq>`l���j�^kF��-��B�uN�<��Tl@��6q3�9��#0��j{��I�a��bd_�2����yU�Ua.�M�JbaOQy�
�ބ�h�0�I�-��;���c~}bDPN��������΢R{��#X���I,d�4����a5y�A���EJG�kkߜ�腬N���f�~P3��Ik�9����y�P���zRp>�3*�x-�
����RX������%j��N҇'�Ç1J7���ٴn�@}%�\���ό�նV'u�,�Wr�M�
j�P���1�mG.�^���(���q��ʥNd�L����-ٮ�^�X�^�mI�zm��#@-9�▎&Dq#�N��{)�~���ʩ!'AQ8F����e�(�J����,�,Â�`H�(�h�H�����@*��-)DᎧ
цS%�ǜv*/�����k֏+6���\�W�±_��>!r.�>O�� @`Qk�Z�����d�c^Ȕ��� ���;4=H�'P�"*�Z�y@'�_�PFtIΑ�@��Q�B��S��6X�^�{��ƺ3S��uj[]����8�//�E�>YMn��f�e	q�j�mg`�f�}��[c�C?���=D�v�"\��T!�u5���|��%�UxJ��*�}�:���j�
��t�@���]Y	�l�O��2W�:��U�L�O���5KIc*�������:ýT�s�1hm��?�R���+�\v(s=������u)�K���󁂘�J�,j)���CX� �~62�1�Q���]���
`{��z�98W��Zm��Vr��zpdc� ���E>�U˝D{h���z9E��2+�xop�ؐ��~Y��M$"W�pb����"c�z9v�#M����eny$��[<��V�3*i#{�i�����B �[�4��r��#JR�/�O~+z��&�i�(��#$+!9��w_�SL,'�X�zX�|���y���+�I���R}vǂ��J��O$,�O�f��7��3"J�!�O)P�����,�m�	r
��4��H
,⣆��3P��s$��@z�0ҞPB�_! �}wM��mi	�T ��C@%y�[˳��;�,f��q�Cޤ�i��?�_n�A�q9�+��^ƈ��d�VTw���8+�^�������N1�=�Zf/?ύ>���lc���=9&�uz�F#ʹ-�%�?	)s�DN%���'>{ʮj^V.�!��Ҁ󼽢��6����Ur�1E��M�U����h�Y��Ͻ�"��p�G�2S�g:2B�N�S�@����F�|a}����:$��Yr��o����;�5#��]�9��:$є�JY,K_DT��K�1�a47U I$�/�gd�d�s�{�F�z��������Z�����
����׸[�iP�=�UZ!N�M�b��t�W��B���
RI�A&'󪙖�Uɡ���ڒ;0�Xn6Fu�9��� ��|5�WY�z3�]��� ���V�=��/�G�!]��43�>G�O�
�6�;&}vd5�W�'��܁�F/yv�����J�hc�n6+�jE}�������׳�*���W��#��,{	�];�&z��z�1�s��-B*�N��������@����s�:�b�����Ye�3J���m���#�r�͙���-հ�V.=24�kzw0�Ƥ�v���i������zy?,��z��u�je���F6B*8&`u����G@���H���^g؇#>72%=�k��ئ�o��ݽ�i~� ���J�,\r4H��ʼad��]�T�_>�*7����|/��������wh�3�ε��,�ubˍ;�>?�9G��}܃e��cr��庂:�jQ�k,�>��Y�l�	E"��c�I
_�fC�KB�������=]��v� ��8�k
�����qp�'���0=�9�6a��wKx�ͭ�9ݔ��v�0�Q~q���p�?�᱂O:�b �I`s�/Y����r#l�◉��n_Ϸ��\b1�I�|
yn|ʭh�<�H���)����/Ǡ���'Cf!I�>eFm���Bٓt�e(��/@Rᾤ��l���A���� ����b2sX��5k��ߓK������Ǽ�M2ݻ�1�g���A�<�@P˞H�����s��ȅ�3ʵB�q?k�V6U�gW�
��*=�@{2Qgw����yO��|��6&��Se}�Pd���OpmX��joL��q7���gSV�pWƺ�'O	R+����|jl�nԟ��鄝��yB�-�g�m���V8#��wRSOq�|�Z�Ά:`�Y@4p����o�!%J�B:`� �V�f�	�so�w� �e�ۤa3j�)/����s,Wӗw[��I����l�_Ff,Y{���K�����d�m������I�(�N!���4f�Y��,y �4�
oXY���A�e�����3�ʖt�ĳ�d}�J�Z�u˩�t�l���C��A4�Zդf��9Lܚs�{�u�S��B��9H^0@��x��J_����IeOF܃E'�gc���Tf���[�ceL�dKm�|Z���o�|�Qt��&$'�m~V��������ɧ�(��/�s����3|[ύa#���ؙ7.Sռ಴�&TvA&+�?CW��QnVT|�'��|�<!c�pc��..<���_�\���|̳Rr�R��h4��\��/�����KMf�,o˽a�g�}w�/�ĀL��҂��`pb��/BS`VXcU.:����aIwb%��E�����4�\.�;� ^E@]p��Q��je�\��-�m#O�٬��4�9;�?|-����	��t$����B�s�%�3h�)�!���7����m�F9ȧ���϶�,R=�+s����ⓝ�����,)�e:�t't\�+���4D��2�c? LOr/����gEW��'�6�
��Nm3��GR��ӓM���#t!�������&�_�'cn���{��1"*�Ya����~��0�=^;N��E�q5��-,�/;��3���ϑU\����ԓ�����]���Es�`_���m7���m)�FZ����:���O�ʱ���"�5�;��^Ñ�kU�����-Z�P6]�U񏳐ԅ�);qP7n'�Ly�^2�U�Ď���w3�}�՝����X+Q۲&�#��
�L1��v�v]ǳ� ��X`	'k�g�_���`�S3�cK�Du)gb���dT���挜��s�d����4p|��lL��"�T��̤8�(c#{�w*5��yX�;���*���)ҭ�./��r	�J�r=�wq�Y�_�; �Q���I�MF��3�֧�����||͸6�Uyl��y���t��Y� �rcU��h�V��C��#7�r���ܻ�v��WƹbF�,w�k�����t����"����Y(�,ț�Tt�p���z!;����%�$�/Yg5�DB��xī�AUv؝��?��M#;8S�rXZ��43��)Ѽ隠��f�;$��!�&��7�b+I�^i���]���=Ʉd@t����A�K�E�p��	t����q:�3��-�^ld�~���]��Ě+r�#\�Ǧv�ω��m�bL� 43�$��Ngi�&�=���]goX��]R��l�o�-�!�p��dd����f�f��۪<�ቸ$�0=�.HU� �<�o���_�5Q�яk��1T���s���RՄVQ)����J<����3[�E+�1��=�l	��k���jШ���I>�.\�a�t3�4�Z@֦
O����jZ,�������:4��E.�
��c5�v��>[� H�zN�HeN��B�U��J�o���7T�~q�p���L?o����Xt�����J�J���`��s���
��u��\b,��t++�e�y��u\\�}�ҍ�;0i&-KyPe��哗9(��DL�g�����ݘ�%jӂs���'�$��^���gU��}��3s�OS#W�uQ��HL�X<��u㤫�#@>�fݙԔ}{�t��O
߿�����_��0��>;� w�O�2�bN����\T_�XR6?���F�� �"��x��U�*G�c�]JT�aޘ�U�|�Ij�{�`D�ڹֺޱH�Oe�;|<��y���a��������~����bA΢�T�00��F[�֣��-k�#�;),}V������7�ǖˉ�r�cd�~Ϫ�g7�}p�8sD&��ȏ�pP%���j��mr�+��!|�ڠ w�`�˯��*3�a5��\Z��"�KvuB���`�V5�	w!�1q�E���C���v�7��Hl�����T�1��@&��v�"�]����h�1r�H�]��1���OkƋ���S1e�;u���?�C/"ίMx-��j�Ew���p����C�\.LC%�0�h��y,��7�~��4��K��AIPA����l�2Cꀙk�7��C��H�&n�����dE[gSQ���ጶ.!�i}Rd}烲(J{%*�M�j�7�u,繇�`�W�[�T�4j6��R���ך"T�rD@��bF/�^:k����N��ෑ�Mk��b&jŊK��a\���&mx&yֻ�O��R�4d[f�%�3W�G+������6;}S:�9(-��\?���.�g�$(���}�/2�pgz��'^����\��do���F���Vx�@�-�#�'z�_1�#��d�A%���s�����4��gM��Dƴ��zC��uo���?�H�[0��,�ڡ�]���|2��y��Y�T���cͰ�v
#44<*��bz�[x�w��QQ��K|7�sL���@9HJ�>���Ѷח�z��F�"|Z@;@��O?������hk��槆k�D͹�k�ҬmC��H��y<�� �Z��>�-�@N}�2��b�̥T��n`�ъֳ�.2�~T`Fz���ɯ���$�-X���ؑc�_s��Ɉ�jl�{��0@�m.�0��F����@VM���	�;��O�o;�R��fC�T(Y�N�+�����;̈� i�g6�'z���_�uhTL��G��x�ef׶�Lv)��8rQ; [��w\�{�Xf��O<�����`(,��P4�Wk+����&[+� "�I��+�tq�@f���=�������o�^îSrno�\�5}??9�*z/퓂.)�n�LB�
t�W ��(��P��ؓ3�/ӣI��ݹJeM�u2;�����ZJ��ȣ�%i;k�e1d��Ҟ�0�5H~="7�[���҈P�g�1�!R V�.ڛ�<3� ���D#�k}V�3��7�d�C���E8��wS ��x�q�=����#�D�����â�G��20VX簦N��=�=9Q1퉫;��ܟ�d����&��;$�%/�U���:"y,J������f�/D4 7$:�G�Ƅ���Q8v��}~,�@�I�؝d�g&(FHq6�A\ی�֮M�_Ƀ٣xV`�mz|��
*߭� �`��M������i�!Qj�����Ύ�<a!}g7�N�N��=���F�E�{�M�i����;d�Q���w
�Gjjzc�Dj{��l��D����K�6�T��J�%�\�(��ؔ�L�2�r~Z���	�:y5�F��Trn�梦>Xb%ፌA�5v��fo�u��K-�����qWD�W^1p�:�ˠ$'n�_%�甧y��+?�bx�y�����؛����$yxk�3��d��@[%�Q��,��_�X�-%r�+$�㚅i
���SY· ��f�g��x<T�F�|�A�{�Z���6�U���֤�;<�r~�0����+Dq�t"�c4K�[�'[����c����bK����3i*ܦ}�)j�}H�zg�P%@I=TG4�&�_�]���Y�m�i���~(�8<`��b��@/���
�Q����k�Ʃ��a#9��v�����j��x�큨B��.t(��S�o՝���A����O�&��
��^V�*�5����U-�&\Yy��qn�6���y��-T��j��&RѲ@�I/�
�`�����ΐ�t�D&�Df��{|B�Li�^��#�Lv1��8T��p����}�?��nn�O����U��8"�9��7��5�1�F}�_��ϴ���:{
�3��j��Y�Jg!�j�xN��<&d��z ;�Hv��Zu+7u�+����s�
I�@�TRN��i�lAH��vJ����<��X� >��X��t��>}��M<r����i}�����p�����9��	����/����M~�Å��L��gcP9��$�VZ4S]��aU�z��{��md��%�	�0�Ǜ��O.�t"�eM������OwꪖU2o:��G�Y�l�&j 1��B͓�H(Ұ��-�_�8XjE��W�s�:\�RAc�D��R�|ro��O�"�+��d���(�m0�nH@@�e�����s���f�C�EX�-b��$�2�kd�7`�� �aN����nD`�=�0j��_gLH^�m��Xm~��8����f�V��s�]C$�����۲b���~�q�Z=���T��>Ţg�A�/K-L0{t����}hO"o�P���Ɛ~ϝ��Yd��IsI��b��ew$gb㈴V�Y�y�@�$�;C)0�Ќ_q��N�h�"��?j�������}���Ǟ�S�9uX��X��wu`�1�n�7��5,-����2!N��q�Y��ʠ�D���N��1:�;��������}�I�6���^�\��B�`�T(tx�-�=�s�aa*/r����.� ��1ɜm��6GVU�bׂ�<Ĩ? E)�G(��[��K�;��?�>� [`�o6�U���̨���/]uߊ�/½��FA�P�N$�x�w�Cqv�VN�5ړnX�1�ëW��}>��l}:(���i���P��/wا��gjg5��ʛ����F�I��D��ԯ|���X��1hĆJ�,���!��O�p�M`����%,�^.l�C��F��0�|#���G��3�i$o��D�}W��I��κ��=�u�3��BU�.�n��5g�YY Y���f���]<�9�' ��5w��\��m]kר��f}��A����ej����A� �� ����k��d�0LJ�r91=�|q�=Ŷ��8�I �w�'P_������a:;4=�f�~�v�(.�B��W�ĭ*h
�qǝ��A�����K�m0db�}�ݮpPl�&v5i���˿v]�׼ 8���I��ph�Ɣ0\�:Ekw릣�b	�Uz�_�'���H�X�ʰ����p2����d[�*N��}~\+ZEț��<����l �7֜�W/���[�]�C߻9h��>��{��կHd���!���K�+�����K[P�(��� �:�fe�\�L�#�>�� Q
[���� ,�R]*�p��K)�l;� dx�Q�Mp=?�H�T�{띦=�A����:Fvu�(0@�MA�ʹi�,�a);oٔ�F��ZږM��ŬxM�S���>o�y m~��J�uܜ���b�t �88V")��}��հ62i�,�UEf���5aC�����d�xA0LO[۰�A@�,,���s��m���d�4,���3q��)���C����V1:�M��6�G�%�*]�P���1 _76zt!W�7�|�o�R?���<j}�s��>DcxOd3��I'1,���HM��H@�L	g*J�������A�Ұv�롯Q��C��x'[�.k��&Q�ۛ*{�����(b/Q��$�.ݑ���lv!yCO�pc��'���z?�O���Z�lDs9���]y��g���Z�D���&��j�`/\�p�<8�5��r�t��ύH��0��y__���񴖬}Yd�,���!�jW���K�}����!I�DQ�~"X7z*�g�Z�Z�bӕ��/��r��"���;���^]����?H�I���ٵ�i_���Z�/]��)�5F� �ii��CE����b��P|B�<�.(M8��+�G���Ǯy�!/4��Z��~+x0�5�+ԝ�,�6�~w���B�$A���n�/�?�T��GA�#����Fc�qѢk!�"{�'��N?�Fʵ ����7�:J!c�WFZs���"��C$����_�A��<�xj�縚����T�~;��ĉȔ��<	&׵�*�y1X���}���r#��St��,��/R.���b�bz��Y���	J��5V�0T?�.�,�����^��Z	6�ݼ��9� �
AA�� ��bU��<9υՙ��`��P�2���"�2�G��Uu�#�
���:�_OUj�r��]�{Oą�ҳ��,%�i��l0���[�'w.�p���c~i&��@��a���/u�ڼU�b�(w����c�G�-�A<�7�v��.��ڑ>�����\����O�4N;E�?yŴ?w�����u+m)G0Ǟr��ʐ���tP~���;Q��I����#zD [�zp�ȄF��IF��T�h��jp��\?�k�l}B%�*�Z�Cj��Y�>��1�Z�Ϫ%,d��G���ɶ��Ӥ��-Pi�;��[��w�
eHѯ�b���3@�HF��i�0��Nff����U�����O����Ó]ըأB��1y�|KT�}�r�p�������S��<�=�7��57Szx"��ilP&hꪲ�"�.-H��]y���].mW�A
����#�l�G�垾5k�F/
zlʆsU�K�_u�b�����ư�U���L��NK�!v��r�M{A��^-��P׹@�OP�Љ2�#b�O@�����T���P��	LF�}1Ҏ��I�A��ɧMi���$h��T���JcU2T�jX�D�f�\�M%X�H5�������1�Ҙc�"D���7�B��=n����F�NO��h���*�w��r1����~n�Q� �����U��?���|W�>ה��i����m�Q�
�a�i�/��#<c��t'�W���A�pZ���XN����X�G�T~[.�d}�����=�"`� ���Gy�v8])G8���L;�=�s���J^�-�U��Q�6K�4 Fc;�&62
N;м���qF2-�3�֖L�JYe���15����&[�o�	���~��Y	�6��f�b�j򩼐`nI�>M,�1�
8��j٘��9{
��'[��{뛉�QU?i%�����\kh��F6��A��'ƹ�=�̊��D��7`J���钯mVT]�ϊ���H+h�<8�5�D��(J��i`uN;�QT'BA�k5�0��`���[dg�N�S\�'t7q[.�|X]$�zJ M�`�6�0��1��"Nֆ�}���'��{Kun#2����x��,�&%���U&G'R�l��a�K�6ߦ~%�]����b�E��S��9����K$�d2�F7��zY�ȤD�Y9)�9��Vn��n^�VQ������n�*�c(��/>�5��K7��%0��	�>c��N�F��(�=�D )!��h-���*}��)=�� I��I�
`�&jVf�U���4�{A��NS�7%q����z4p�1�P
�d�${��	�I�����ߨ�����{e��XgSE���X���� ޢ���J���0e[mZ�W�
�l���߷5�ĺ�D�A�pzc��\c���!�gF��p�Ⳑ���6{+}pf=��u�g��C�lZ��^nꥨ��*Gkɉ�(�|>�i�lt��?��K�������wi�s�`��C��<�<�/�p��J�!�N�/[���H �*,V��1�E��+�T* ��q��g�8�-�%��%Ԛ{�/'pD��
��죲���Ȋ����;mծa������{��f���r�O��?�����1ΟOmҰ!����b9(��� �A��n}�Da���}D'� �LH ��ї��4��vП��=q�vq��b�+����	�A��Ϊ������<�sw��҉���l7
�%Jܘ�!��֑��It��$؊�Y��V����5�M����E$Z����+�A>�m�[d�M���ָ��
�^�
��ޱ�A��#�A�@�X����*5�v�0�ʟ��琨�@�4�$3��mf�������σXG5���ɇ�,�6{=3���@r�˞5j���u�-�j�3��F��۲���A5���ɩ�5�	�=qo��#qv`#Z�p\��� �ծ�[��b�gQҽ�������UE�'Gv��������JKެcH�:�>϶AE�e��݆I���-�����L�n���������,xW�q�e*�&W}줅;����
|VWxZZذ2��"?��_O����$2�D��d��э�z�pOE9lZT���W.���
o1_�ȪU�0s��`l4D��߮Hbl�oh_<v�����:]�j���S��r?�TA��6�8	@��8�'�D�/��ƐD��ՂAQC�<�gM��l�} �`o��`[/�,ÚeA���eop��Q�/#�B՝��Bq5����7Ջ��SlJZ��W��^�����r�D�]�$���!����{*�3й� H�i�GV�U�	֊#ݑT��H{0F�Z.W`�K�
Y�����7ݐB<?����d;[w�?��l�����#��P����<!����S�eox��Xp	WܣS��Ku�mdQ�2C��|����L���ӫH�MF�#C��k����:�ܐ_�F�uX�K,����;�9��#x���h�[���>� �W�Zs+�^z�w5��ȖC�U*�d۠^�$�,�B��]T� �B���;��)�.��藾���oK�'l�(����zQ?�3�_s�g���Eq��R�-x�Ά��.�v�x#6L��1v=&a$� ,�j1%a6g��>���2�j���>8�N��jI�����Ldo�'��� �?Wg�~�����r ����߹h�v�\�ɇ�c5�+�����~d���;3��x�%���Ӹ�����mL�x����c%̈��A��U�0������@�K��y<�jUǞ�_B@��x w�r�S-9`H"�-b	 �}�"�j�t��Hn�=���ɯ��AM|Ӄ8��%�Ċ~�,DYD��	i2��߂#X���#Ur��I�!�W��
�
'�֮�͚�ۊ���>�P���a� l�%V��'��&��C��V�^꼣�=JS�__�u������cm����2������x�(t���ڞ7O%qz#Xu[�@3�6g�g*�`�J+B`�~$�����?�}Ex	.U$`�=C�m��qP0uV�w�����q��Xe��F_�i�@�c�֣e>�_�RxkbV-����@
6~c��b2\{fN�d%�Df,ܦ ni�չ�a�����t�t��m��?�ФhȆ0�&�[	��P��lR�Ł�s=�xu�Q?�ڗX�B�Y����M����pb�K��V���h��)�>q����� j$֘��`G������q����<ɐ,ӑ&��=o�u8���,Yd�@$Qi嗡�"-�!��1ě���)i�H.nc=`U�F�i.
��0f�7D�
l�F1��2������ʤ��o1-��;���BY:P�#���a�� ��0��?�	�! K�=X��9�[M�b���#�y1�m�5��)g�4�-N�s�i����.=z�����2��A�� f�����Z"�HjH����f��뎸Ջ�:�i~�r�Em�U�u�'�	�4fP�g�b3?��`"T�
�R��֭Y���`͌j7�7��KrЭ �&��3�������͢���8�4�?73%ǻU�1�ѽb���1C�?�Tf�|��OA��UĈm����j�� on�yL������Rkޝ� �r�E����غ��]�b�H&� �W����飶}'|�s�B�w�c� o�'�w����҃e<�6m��b�;R��� �Noݤ���Wz�S��k���L�3��
2�r�7�fѫ.4��I6���&_��p�����zL��"d#��~P9��L���,n|�pc��ײ�b�u�B~z��;������C�9��7�R�7{�f[��|�a�����M��Z>-�����*��lDE�s/X��'��������B.�|�}�̋�H>�[���mF�= 6�O��QX�m�����Ht\��{�͒�0CǙ�zDi���1��+D`&`>76(��;;b�EU��������Ŗ�tՄ���f������J��������k�q�����8Q� ��hAq�idqQu��p�#��֚k�{�(���T-Y55���)S������u�d���/�H
0(�����8��
}��:���'�@�����;���E1�P��{��h���q�7yZ�+#�`���E��+ǫ���W�Wlo[T�8
^c�	.D��/(��F,ӎ%R�e�Z8�"�|�DA�$}�(��!8� �D�~[;wI���)ٓ�$?8�A#��@�P�`g�6�a�3�5F��7�9����E#P���*�B^64dܪ�����v��#7g-f"n[;�M��LL|��	;�yRHŒ��b����lb�ғs�#�}J#4!�P{������W�'��iQ�Z�����\��"�O��ƺ�m�#�!�$�$P.�4�R
��49����;�0�)K��,(�~�Z-�<�%�V$+���H{�^�|u[��>�-=/��C6D6��-���ݳYq��ڿ�X@�� D�&����W�M��Z+z+�D4Tq����ag�Ai۔T���?�p��t@���ؘ�BW��8�'w��Mư������n,��I3��{�~WP��l~��m�`ĸ�G�r�>!<R�l	�m̈́�C�ǉ�I��p	�Qϋ������o��u������\�#��{�k��jZ�|/�M/S��P)�FB��
���k�~��`��|sȽ�n9�UY8p�oQ�q�l9H��_�xpY��Tld���g��j��Z�ũ�\�&8n�R��:�B�(�Sq7N�äm$�׳zf+(�q�8O��8,b�4�����h�m�7��~���GG- [h�9��^��Et+��7�<<l��:���+��eVE)Zz�L�4�����h'���/e11�k�/π^&��
}���?Co���.8�!���I�t�@L�$?�Z9�&����j��dkp��9na��X��w*7���5D)�0�<`�6S,tu��e����"��'}�)��>N�颿�,ߔrY���M��=�8d�c�D�p�H�+��dp��l�P�"o¡[��3a(B}`G�������+���t<2oŔp�o~ty�����>|G��������q��
Y�Ƞ���-���E�.�L`vX���<��9AR+b�ͤ՚�MA��(�gKJU�]���Q��M�,�1J��9��P�ߘl�A�����;<��aݞ�.�U�f.��O_����Q���8�"��}/~�),Y��|NX��}�� �<��c��?���z��2��x%^⃡{���"3�0�r\-/6�z�k�@���-ЙmȡfJQ�*�5�Lr�;|�����<�ŉѴ�D�ڧ8G�0��_�:c���WJI���i<�����=�I��}T��)�o *��E�D�l������ �Q�5�Xo���!ʈ��Cj���E�\���Ӓ�J#���s�U2+�h���V�q�M��a���� YZo�yъOo�������ѽH��O��du4�fyrecs��:�P�ԙ,�K!T�5�(��ZV|l�Ɯ8��6��H�(�B���rK�̓J�[Bgs�C�J��f���#���_j�F� g�}�A�6��&�U�ʡ����Q-|���W��y�&����S�({��4H�ά���s~A�̟D^��ƲudG7���G,s���УQ� {�74�D�����������E��4��է�z���6�DZL�%�MWD-�l�A	����L��]1%���3D��e@Z���Uk\ qW$6���
����w���Y�پoMK�O���uvb[Aۨ�P%ww)D*Y�yՌi��>�ą�W�*o��Z��\��vO@��"��t��	8�:蘜�D]��7�o����WQcnxmML�k�4�1�S%�]��(���%W�$�����VV6���X��(�1�_=����pJ�-���FN>^"�X�-64p��o���7O� ���Jr�!Ȟ�����/�)S��!,���Q	��ɤ�V�!�c�R���l�b�Ͻ�\���Y��w�w�GH.��W�뢮���Vb`�ٕ}��X�ۃ���KM�j�Ր��$8��L��~��9�IZ��^S"6]u���&�:���_2��I��5�
��*�+��2�q����-��i`�VS.��X��!dƇ_�9�Rɉ�%�ϛ�H�{�ب;��P����ʉ㉁�a�i��u&�����;�%��~a�+^��Lk�[��iw4+����ҭ�Sh�2oX||����F�I�چ�	T�kMt��Y��6Rq�U���ױ�����h���d����I�䣖��M�W=d��pEsQY���)Z z�>{�����q�[c�&k��;��QE�i5�˜K��8mS�~�EUȕ�kB��/X����L>,�v7�N���&Cyj���B��3�?�Ę�h����\�x�q>��[��[}QM��'�F�y��j�~ZF�iv}E_R�
*ը���z2=|�$�O���H=ݼ�@I�:�n�A�������* B����H.Im$_Kw�{�� �2%��!����
�Yq�.����"��ep6�+���dk�I��>|i�*�d9�UV��eZ�_Y��qy������^��ݼX��<ai������
��jg%E�L����#�<k啑��_D[r}ho-L8p.�1�g�_�;�B9a��bE��X._ eޓ�Z���!?�܀)�������c��v�9���+��^*[4��S-Uc��~RX2������X.�H(�I�����)*��--ǴeYW�>��;�RԺH����*�ތՑ:$Wx��
�L�o�$���ucn���F1h�?@M� �DR�
xik����3���΋� �:��}<�o�#c�or+����}�N	��Ĳ��{3�,�)�����fM�9�b����^�Lt9Q��A��Am�C&�4e�z_�D�t��s3�EݮkFAg̗�D���8�h��G�U�c�i^E��9�����][`�������2�v�K�.�8d�Qxbk*z� ���'����E�e���e҅$w�a��59ލ���~d2�s�ҐrL�ǪJH�Dx�pz����������
.*��Id+��=+���ܼ����G�5w��ϮsRk�V����.�궚�!%^�uq*:��L3�����;TW��������,In���=���k�txD��3�`'������[؜\��rvtL�kI�g����s������b�e��F�w��φ��7�_v�E͝�;e�=��Sp�Spv��PrU1
;�Ӷǩ��?�/y�Tf8_���N�Gb�S]|��b��F))w��`�\y��׬X�S<�YwC|��wRd��HO�I�;��{��ـke�m��EL<,��N�!p� �aʄF+�&��9U'��y�����i�m]G)S�M5Y���["���+wC�V�ڗ���t(�!4{2���x@�D��Y�,�vP�?�0WL�kn8��������=߸�=,a�!~Ƽ7��/*�؟����nX*};��"���I@�>���<[c�p��'ȋ�	 1�3����Ҝ%Gc+�(9��<06:�$���Y��7VU[����b�o�0��V#n3
Zu�d�$|N )��C�,�<(�΢:���s��r�Z,���ќ�>����Y�B�`�A�B\�gv�@���"n�l�Ł���;��;�e$��e���u���&/^�w��Kj��88�M�I�w�`wD硹4��Z�]��M�[ ����Xp�	�>�Q��OEko^�9�&x&^LkuSJI`���ݼ-]:�iuӢ���k�I+���M[K�h�	��f�ho����[�K$�=�%�fK�@ճ7�N(�ϕ,tW!w�8"ϒ�����>�Va8!�W
5����ҁD��e�$%�^�w��;�Jt��Hᇌ~~@��w�_��w/b�*,�X}24c�7"�Դ��ɸ��"�h��Y�ÐxM��1���J*2u�״6@g� ��������^!�E��}������|b?�iV���^H���N�G���WBן�`6h�����$���N���Q�����1iq��V;��f�5f_����i��G�4<�~����_I#����!��ږ{����yu2L�A�J ��q�+`�� ���SP�����G�a*�	�Q3��h�a�փ�p�I���} OI���W�[E9x'?=�=�"X�&C�KH,�aX�;�=���F�a8��\=M�P�8��i��6f��U�ټ\��d�p��b4��8H����L��N�����pTt�b���P��
�6��w��m3����t&Ȥ?x4�g�]�5L��Y4��C����� �N��x�ۆ�;'�v� C�ģd�������Zw��6��gCA��`�kiNw��b��9��U� ��
I���0����A%�)���.hs��TL��6�d�ɽ���t�`�Ix,�"V�;��F���.��o�����N�fqb���a�g�X�[�!P�8�C��u[�$�*�4lir�$S�I(����*�_�e���a���=�����u�B2~��Ò;�Ax����OU"�>!�DDVh��6����d�ʐ/QZ�I����J`���k��F}	u<�G�v��r[L�"����N�%(�nv%�2��I^�Y�ϘB����y����; 5��]�i�5v/�kxO�@�)���
�����H*M�#�
g��!�EӋ����A��_��X��x�:�	(�ǜ�l��VF� ��(���w�aB��-�����C���<�"8~rb]�;�c�hx��ӊ�A}{��1a��=ڙ��F?̽x�3�#���{ [�x�'�ZsMc6��]I
ADܱ������)%t�[�8���
�4�2JL�&*8�rY\~�$�>�e��1�H7���:�K�xr,��TM�#C�F�8��F(��g�/���
�(#x=tΗd�[a�����w\\R�/�+:��m��������fI)&)Cr��O<r����#U\n�JƂm�d�@sD��P�!ñ�o�:�M.��bu�(zk}�&ܺ=K�7��&B��E�]��A��YJj�����Ha�[��ǒ1�2�??���-�Z�P��n�EZMD�nC���g`X	��%N�����i�R��?�`�$I��^](���nV�l�N��� a��y�iF�h��h�Z8䐙�?�k�����UØ
�hٿ\+��"a������E�հo�6sHac� ^{O��C�&���tF@F�.aY@.���lx���e!xō��2�#�p=3�4	�N}ѫ�ĩ��2޻]����Q��%a�K9v.�u�@�]�eѵ^Ԓ^�W/�3���K�e�����6�kB���j}Sx�?h�aa����u�7��^5$�b�P"K�*��� ����5�VV������Լ�vPDS>�!���J}�u���kl ����B���.�y8��.�g�ԏ��H/���6e���w��)���H!t+Q��i��]	՝�ʣề��޽b'�x�i�_F��QƤ��̯Hh1�A!]��|�V�o/�Z�*��|*�Pn����.η]�I�����K�o�r���b�y�Q�y�~�q	ׁ�%޳
I~���	Z���*���� �X�R�K��n{� �x8����9�g&��SC�����T����6�{mӹ���s/@�h��j~�V�q�ABRP�R-l�ă���|2%X�<?Q"���� i�\R�M�]i�(���j<�m���@tBZɺ4�OI�����y���ox{ۙD�y6fd1Tr42�>CC��A~m���Y5K�>�Dd��[��4v�O�Ћ'
h�#%��{�_B�,W;����fk��Կ+)��= ���fmZس(O�N̞.�s�B�x��b��Ъ̕΋Mű|g�2h� ���}P�ac��.&)��'�4���H^V,vuNpu��+��Xk�P�#Ъnu��6���G��Y�{��R��f
	D��CE7!t��]�����y���Z�/��W�nKa��,X�k��.����i�t�J.5��7��z�߾ҙW �ʡE�黬��@���".k�&������6�ߜZ�+/|�4mW�o���F��<������!	��0K2F�:'�<@}j�-6k�tK�<�aaP7W�k;%I���?���\TQ�tܐ�t�c����LpN�a8mC/6����Va,:��)�F�8�Y����*�Q��%��s��n+z�p���?k�r��6�a!����,/[��r��m�#2�+�YtG�L��|��@��h�R8�@�c��\V&�sƢTq�{�gz-/#�oJ�Y�ڔ�{��{�]
/�z�w�vҠ����+�;��<�ܳ޵�)Y�h��ؒ��"G�I~��@n qb��,�״�lQn��]bDo��H6��IŃ�]_@/%��$r %Cs�Os��J��OQ�"�����M�����Ct��m���,@#��{
�� ��GH��������.۝���nU���S@����§'x޶c������ն������1�e�Pe�5�C1�A:����u�X�?p�3����=��ҙ
���2���ie�;��4���[e+��oS��g*��#}+�L����"G����]�F�8����;�
9]�jH�)�x�&�V�(�?���y��;����*�ym����1� 6�o|
��²�%�����򵺊2�rU ��k��؄#�3��J�OĲq�� ��h�f��G���Y_Q�d�4�H��`p�LZNf���K��#���n�8:{jν)jE�_R���}Ն��p�E�#&%I6�ᇁl�U9 �ʠ����̊H>�,34�~��r�WhA��R�G��p�rn i�y5�˃-�xY���v5�2�b�����x�����|1w��~�X�Iƣ���HY7vNL9����:������,TϘ'�0v�J�l�_a��%��X3��C6JK�~󫹸�'%q�N�uH3v�+t�v����&9��	,@6	^9=�0��Q�WT[IH�W;���#f#>3�FI�M�o?[F�E��P,�Dm��a䩧� ��5&�ګ�رB�P�Խ*��.�N��7�8{��G׍<�� �t#wn7�,Q�W�x���gG��!O�J���t7v*>��(|$��"L�u��K-~�y��f�Y'��q�k�}H�n3��\K�1�f�������]��S����h��h�:w�t��m~�����2斨)���A�任k)!�ְcy/`c%�"T��x��䄯rLk7�\�?Ey	�՜=Ö~K�;�[F`a�?�-������胉?k���ʹ߈䑳l	�+C$oa�!�?�{�q���Υ��ƅ�l	�_�Ǉ������p�ʬ#^1�D�Q*y��V5J����uq�x~�(��y�9���3t��d>N������$z�w2 P\XU�K>O0���&6�1�2�^�#�M���3�5�NL�p�XV@}�[��?0��^� �����?;��`QR���"{6|N��0�.�qfY:?:���$�*y!�]��툦�]	v����ϭ�F��(��h�e1睉�(r�@d����_�e�$Z�i�rh�KF	9�r��i#{�X�U#B���"JZ1uV���	�4�W���j��u�7����)��?/�8��.�"|���������/>FRuƏ]ko�&p�L�����!���7}�1	�*���?I��v�Υ�.)fd���k���R
�*�|sa�K�	`=�	�P\�#������/Z��tA�`���Ie{�4��,w<)��̉�g�)\�E?k���2zw�%����zTlu,R���#�z�?��ò���ƋP ��~�9��0x��KS��(;��!7������/�Z�í �^�t7%Htԭ�
9PH>�@�7ma��@���\��ΈU�4.�Ye�i1Y��߃B����p�.S�ĉ'��2���gL��|�M@����t��U����?ʐs�-�t��8���y���C��Ԃ��L$J���{�R�|�����G�9�2��-��d3�}�Qa�����XFU��Y��1;ۑ����ⶡb"�E��MQEm�mD+�Z �$=��Ŀ����etۋ�e�^_A�S�p��T�Be���WՊ�����{�=�;�
������C'�ܩ�i�6Ovbe��:���G[������|���T�m\�gsi�\q��o��	Q~�Je�Y��'���5�7ր�%iԔ��B\n�����	WW��:r�p���������%ﮧ��V[��s��ꤤ����m�7��4�ҾM���cQ�w�CKH"�ػ�#�$0(���S�kiq�E�W 
�Q�e7/��ǒ]C��i��w�M��(��JFo�*=��'�'*��24<%Q�����G���UNYg�d���P��0N�]�s;͹���6���d,"Zh��D�ş��3��i~��Q��'�H�䱬'|\	�j>�D���N�wA�C��P3�q-�Y�/�j4�5����C�W�,����nN��?��,��#�+^���":+Ap�,����~�T�NF�R2/���hUl�r~�o�	����u\o��HaHr _4p��%��@c���*y��o��C���"\�;Q�[c�t��ؖ���}#b��v|1���Z���f��%}�Q���:�2��VJ��i�v�0�ZNyETc�V�4�KN!��{ْ�%�_\��.�� ^��nZ� �ʜ����;�؟4�}i��̅7��?WR]���ǜ8�����-"1[fjKt �t���5�7�F��
�1����iՎ�=��g�+�8�Ո1
�4A�Gp��n�HN�z�2^�P�{��IeO]��Ols O��]n(k���dIF��B�����б�������'{� A��vr树(.���	/�$�,�r�Q����_�U�<�4ߤF3$�b9>z ���_&�3������Ώn���r�Fպ�8*dp�-x5�L��'� �A��qFl��՟i݄�}�ͥm�9v�9h[x��G<�Þ�a%W�Ix�sk���5ݸ!F��BW��V ��.2窱>��k�@u�������R�N�<*	�������F�R�������8/(�1�:�^n���� ��2����.����W/ǎy6Ѩ���� tVB)�n]Z��4������0�"e��x��V皮<>_L=���rA����`��Q�A�J=ٌVӤ�Y���T�� z�;w�%U�ϟ�oP�� 3��d[�6h~0>�Pp����c�O��K!����53�䧋������C�At�$�Ỡ0�i��m���m]���z(�,(���:E�S5�� �,Y&t��az�B�2Q ��B�b��#��9pn���-���q��
���Q�n9�MK�"����2����Cw�40u���P}�� Ͳ���)2m��bHu�
.*�N����r��:����P�y(�����|+���0c�&�w���C%[���zpC���7�S7҈AE,��AO���Jc�XbA4���E�}��|�IT���Sk�T^T�L2���Gq�L	���B��
7T�zK9���8E�om��6L�{��:�������������ܤ'(��;��쓤Vէ�hj�<��A<(��rX���!aa��)��F+���t��б���X�Β`M��H�ޠ+thӼ 
^,z�����X%�.�ֻ�:e�1���#!|μ�e�/{i�e=S"r쟴6��"�c��a�Q�V����m�����s�T�'���s0���0�_	��A��Y�~�`�F�\#Խ/���i����?ჴ6�fW��o]�7���0��R�p�jhx�Fx{r�U�SB��:?|a1�"��0)]�a�)��9f���<�ǘK7
u9�~u�?E�G�D���cjH�oyT����}"�Q������^�����S��IVèI1O���� Q�g�/P1J�k	j+�-�t��~��;�Q�M��z��E^R!���-�u��p�E��I9�3w��E��ַS?�c��x�݇�a�Ɯ}0�"-�����N���b�گ��z7N�8�N@8R�O<�H�{A����rK��ۜh���q'�9��J�<4p�p��n���Ѵ�ށ� ��u�u�+X��q��cz`����8M��E�q|�Hv>Ozt-���Rǵ����G���X����1ܳI��U8���p��C��4ԓ�=���M�c�b�dr�I*�%�t]7�Sn�����k^�a�8ʔ��ՙḋ6����XN��G�d�vJ�!w����ǓS��_��U��1)NQH��So_@߃m��/|�pWرƆ~�:*��*�΅V�Zr��=r⺱�C'L������6[ʼ �m�����U�1�q����yI�-���(7p~��9�,�Ω���e��L�S.薴�m&d��+Χ��J��p��?��o�a`��:��l�f��*�hh�g����w��,f	'�)� ��>��Tee���ٶ>t;����f�}��7�:U��7~d/���dlm��u�A��[�\]�!���]-c�.0l���jV��y	!^t��|g�h\���=��cUqgLP������[.����M��T���QI��OʠNA[uS�#��Y�[�wjh�[�x�s&bfe��<���´UM���ſh"�\���Uܰ��_������-Xekõe���z� L���nǲly��l�+U��@m?AW6�3.ģ`G.�e�i������?r���1߃�~�6�p�h� �T�B�ѽ4@)���Z�P�HB4x�B�T�z��˽mf���0?�_����c
=D��ך�b�˳�`����T�~��2΍'a[_'�`�"�r+�M� ��sz�@P��$�����>��Mu���f������v�h9JG:#�&���DxU�؏.�Q�e�ph8�I�Px��%��}�/ʲ��H�B65w��z}|XT�I6BL�D�,��N�t�B��}�P����2��^�(�>2U������T��d3���������|�{"p3W��|�/�܄d�#y"�-86?L6�k9p����~"�A��f����i�Rm��\�f쩘�c�3x�@A��}�z'��E�9�h�U��Q�ɛ���Xx�x8�&�Q�/g�]���_��E\��.O�=1~w�Y��6�IZ��lMp�TyU��z����� ��;��G�
�&���/oC\���{H�,��=�\?��rP�	��&��(��V�b�����;�[����;j����q&��'�~�ZG�� Z�a�MUȜ�(Jj�5�ؗ�A;
�R$��ٮ��� sG�2����>@i\`�9}�(�m�����]kx�a;���En��t<�go�цz2)���'���<�a?4�:��u̸%�����#���6L�Ӫ���,�R���4�ǣ�@��,���k����oO�=})�/���x�SN�Α��U���O'9x�׺��C:#���b�q��3�jz�a7c���x$B��{�C�y��ԣ�r��Z�����N$�2���AR�G*�LϏ7V�Ęņ�GJ�������!��wpͮd�(:��d��gpu�����uZ� �me0��&�Pr���}4<��* >K;�;�Q���+�[�֟<��c��r�o
G���
\�5�'�A�52��Ӱ��eV���h�������e�n�2Q��j�د,O�z�t�P���Ğ�T<IT#HLgX��hD��i���~���e<�;ws9�Uŭ�������j��FA�����_$��2b�T �d+Ɠ���
�@x"��p�`�T���J�b+)�O�xq�!�w`#:;̿������d<�\@R-7D�  �#eo*�`���y�M��.��E�����E�%��0�.����f�>��ݏ3'9@�8/^�?u�ս�
��t��p���v�I�F*q�����	�jJK۲Q�l;^���0�9��symY��7���[ͱ�ʯ��G%UuF��RQoٳ���O-݆:[OtErG��X�����5r�����N;�G�䋄7A��"-Vo��j���iP,�e�"B%��֎�|95�t�� 	A&���Zx�ڑ�_���F�u��C�IZz3�<VZ�F���@v9Vt��|x4N��~���h��U�ȼ�YH���������$@�*$�/�R+ѳt��\�(!ab�W8ͅ��|��4����J���.Z �.gIz^���J���݁P£u�A�*U&�L�w�n��j��H^)B}kc��n@�u̝�@�XW��O���!�~w��J�I<d��-E���}�W(�Q����+z'ۏ�v�Ix�&v[]�:u\<!�	ߣ�S�Kq��@�{�)�ɂi��v\�<UK�F՛�Wm��S��N�g�Z7''�X�W�Z��V1{(3 AP��j��� �+����ZHNǼ%G9O��x�Bu�y������zW�Ra�s��2(�	T�d�U�VV`����(�E�&3H�`Nz7�q�g����f��ֆ֠�C�j��Vt�{�}��.� T��ᑱ�nA�׿��3\Bn��xVm�̆_��)�%�>pAQ�&�������G$A��dT��3�V�=�����^0�o
S�VV���8��R�A3�<dN�)�U6.�g�Ey� ��玽��99%��YY݈�o�U���y�"��Ƙ/|�/��W���9u��W΍�܆��	!H���1
��Q�����	i�v�0���S}�+Y��/S��J@�7D_��AL��OkX� k�
f�����Nͪ(RW��j��UX#�?�"BrQ3:P�n�.�+_o�]I�ڨ�I��ٿ�G]�����KQ_-�[݊�q�Xn :I�c��*�}F��r,K�
���2h�ZKǧk(�M����?yq�C��B5ji��m,��*��V��D'��pt5��8X�Y8~B?����O��tvՒ�_@��u��1�5�]�[}�]r��������ȸ���K�Kw�
�~G���1�`����o#U�����s4�$��뷫є����@c��u83I�L}ŔP����+���;�_�oSl�cuX�8�7�[�(A�9��.T��Lg]=5me��U�uO9;C�"��J��˗�qdޘu�G)'K�,�i:�#�X9��o�W��1v2��Lq�b�i�X�e8鴬�O�E0nĜsOKļ�����(��-
���-jׅ,��n�b�tt��;�˒�$�!��T��-�G�����HQI��*��F�P�����o����Vi_��5)uO�ވ6�!@�[������*Ԅ� �'�gF�3Q��K��޺l�t?q�Nk��P��Gpm�3*c�m ��z�/�_��x���vY�Ԡ�����-F�DTc�V)���D���R��Bb��:��+�ǯ��B?������e�D�����d�p�RH� {�����\|p��
؀�QV9?�T�*5r5p"���p.��5=\	C@��I�E&^U|��A���So��c@"	%���^y�+$���	���/�c�t�PD��6`�\Q�yr���{��O�Y4�!Ӳ��g�6�ml2���Y�h��0=�7\�D��{/(��'����+�B,�O���A���GD�XP������]Y�)ԏ�Â&PW�ޱ���^���FΝ�Y���!-0p�$1b�d۾�D�̔��b���D�JB�	W�FR�d��ګC�D���G�X����'nD�QQ�����j>�O�� �3�W���Gv/]��n����Ú�&EN4�Э���g���5k87�FL����p���ş�T���i��!o��ֆ�ߞ�]�\ގl*C ����q�׫{w]��@�l�QK�����|Z1w@��`��N��A��#���q^<c�7^J���q-����;|���7(��ƹ�
;�A�#�M����8��[�u��9��b&�Z��,�T�g�b�)�x��M��si��\�jq��+�㭕^S� E�}W�Qj1D�@ߊ�����&9�����|�
�� _�Y��CZ<x�����A�7s��-<���)c��NA��r��<@QT�����:R6�<aB��z�IB�̤-rj߃8	ES��,��~��ۇ,~�����-ztI�2�.����>-� O#pǒ-�^��rѤ%A���x��q4�b�Sh�;Ї��M��,����ć�fYN�B�!�*��N�����b��w��A%���T�r�
���5W�#v+�Yt�~8A7���y�����IΟ�d�pRRx�������V�os�r��*�cRێ�d	��W��S�D�$ v@�)�K���7IA�{tnlӕ5O�S
�^%t��E0$@�=�[��|2&�询��7�����7=��� XL&|[�����:'� ���ɀ=�jmƻ�{���{�$����>�-74���5F�V8�nz%�d����PTIF����c�YB�=��s_ћL�j�*�6��r�r�q1�@A1Awh�wB�S^�[��ETľتA�;�����{B{S6���M�#	��^��*���������i8kr�g�./�t�-:�=��y�G�tdn�x�y(��H��3L.JB��H���ΎU>��
���jq! ,���A]:�Q�,���^�R�����89�su"f�(�,�$zq��!l1Wd�b6�`�^�2T�Hrc��Sg;rW���u-N�/2�#<btҴt"�V���%�J	�UN����;��)��E�#�z�s^X5�W�ŋ"n7B ���H�]�;u���oq���g���i����ǮqQ�|�$�"ڭ�5deŸW���t+IJꝨ�?��a,���7d�
�״S�qzuw���~�"~y W�=�/r$3�Vh���f���T :�����F�K��ϓ],T�dlk� CM
�T.�c�}�u���z~z~㭾q]d׺�����z3(���l�%<�~�Ӆؽ���g@t�[�-��􌤲�K��&��c����x̀��J��;�]�����Y�^ \<q�p&�&�t@��:w�v�ќ^Ɠ����K�	O��t� #� ��=��9*��p�.4%�E�İ6�o!ݏ�Gh��������i�r1'�7�����45��4��BI��ϋON��>���<He�H�}�7~})N��}���X�M���,T�ϗV�_�t(9��E�a���i���ȴ��� ��0�����Ob�E.8�3�Q�ט�����vO�����~�jc;vv�Ubtd�6(���zh �"n�bK�Χg�l�L����H�.����ƙ�3_b6z�f�Jhހ�Z觙��0����A�W>UMO��%��\��e�%C��5�)��3�)�$�&�.x!���T&�ء2 ~�D�g���J\�~���+����U�\�*�y%���y�2�?����e����@�y]�Jg힫�5����YͲ��9����|`����rۧYg��@O�B�d������:)d�*����u-w?��H!�FY��u�.�ȿ��0�.��ǵ�o�A�o�����W��ap5��g-'FK�Α� u��Eӄ�s] ��ؒ2�E͒����A��_(N�,H������p϶�Ģ��T�-��ɖ+��k�w������J��@\�f��Iw��=JO��Ur�����y�ɱ�s���f�BJ*�G�$�] aS4���~(ZF�7ł��oK"���=�?Q2�SHn�FE'v��h8ۆ��F���iY%� >�"b�)DJSN�����4]��A���K��������5�F�Mϐ�7��:��n@À��3��F����3~ҮG9��V��x�w�/4�`���hy����~�`ʀ>�H����/-_��xC��,m�"d,-ܶS$Q�7,��)�Yt�UCA������T���r�"p�h�Šh��������bb�#w��:������̀"U����ŕ�	Tx��f�`�j#��X$�'&K#���uE�&��ؘn@����n�PEe��O�� NT�Db�M)�0&+�����n��A��U����lX�#���8��}?�Q?�:�m
̊Ke�F�HJ�������Y(��k���d�?"sћs�hQM.)"LV)�$�fᲸ��x�������H/&�n�o�=7��.��Wu��)���yy=m���+�+��tʂT*B�ֻ�^x�I�v����\:/���+b[�0��V3�$�Md�&z����|�?�ڍ��:�A����,�H��UO�ʀhc�/#��rE�!��{��K�5��/�
��-'�Gb�qc�a0�����;&��u.!7����E�A���A}t�cښ򱰩]
6hl.T����|!cP1 �w�`�Kj��(D���A(~5\ۺ't�yt�k����\��z"��E���݋�苷��w~���;��X�����S�u؈�r��ك\b�:_����k��~�h���v ��ڥ,�c�Pܦ�V��@�6���ऑ��a�ת#Q��u��H-�������Jj�Edlj��m/Z�Xe�I�ȕ��[�u\�͙0�aO��W��ƹ҂�b�a`��E�G�=T��k�x��-bȑ&��Z�j�:�R{_'����h8!inܴ�#��N߯h֔�A��<?Y
���y��j�)X�<� *D1�sZ��ݥ�*��ƅ�>���
�Yv�%���Ξ{�gى�W4�~�nQ�Bb6G�ݲ�E�Q9�W�q���s�F�(��^��������G�%��=+�L`މ$����)&�(�$BԻ��)��ܕ���W��W$oB�N�htݨrf�!�������I��]Q�C��et 2$ɓ|�$A��f{b����ܤ3a�c/i~�U;nH��7)� Ƥ�x5��Rx�}�/1�ȴ�P���31'n�f���_��q��S�pJ���">3��T~������=m�z*��>����-ɿ �q�3@�-����;ݝ�l�3���[̏Ng���b�$C~�`��ӥܓ(��vmB�Y���K��^��Rn����_���l�T�7�m�Կΰz��^ ��+E�?�<A|���A�� ���+t��ggM�[m��vc��5�Jȭk�[�#�X-�/i�!b� ُ���>�͊J��ԙ��A.O�ڴK�����6�[�U�nx� B�[ܷ�C6��fs�.��}J �"��j׎��|����o�������%��^2�q�U�9O�[�휔���r�@�kpY�
2��|�X��D�fd�6+��F+�-G>�̹Iw���p����^)~#���(��p���[-����:�k�CKP�֢ b�	<*5�����.�0_?�ߖ��L���N�aiܪb�ӧ��d��(�K��M��$& �i*�ב�����.;b(ޡ�1r�� <]\���z��>�4~Po�r�Ē	�,��N>�`��-��-�P�H�D\lȯ9�K����9
/�X`�:�+O�5ʮq���w2ۆ>c5�����|�nF�cG�=��z=-�8��T�N�y_���S���̍iƀ�ys<��ߧ�/����q{�eg
��B��U��'Z�;�$t
Qq��پ'˯#MTc��{��E�Y�;`B��*�����:H�	�cM[�^V������hk$9�ŏ
�zZ���!�K��DmE���X�xO_͕{�<��]	E�Ι�gV>W����� �%�ӓ��lz���-��d?�ƆE��!1{�/�,��hv�&�?l,����"��N����@��Nǵ�����j���XQ�6�0���VY �%��*�k�:B��ޚ:b%^[������@`�~@׶8=���ko�Du;_�Y���wX����8e�\�`h,u�U��t%��7��_��$�qV�����y�����0�*~�5�B���/�|��r�����S'̌iS��'F�u��["0_�z�M���E^��Z��B�C�އ���8 *��{�ǃ�(�S��9U:��,eܾ�aѺ�E�mp�M�6���"cj3�������/c����X�,��2��)�\��ݟ�؄,��[I�nT`����
�ӆID,40��I�*mEE<��z@��j�{����U(��. �Sa�l卵{���+���הH`� ��T�Iߺ�܆��2�4�8ܪ�O��&ZA�����c/�^�����ځ�qԕjC��/�A	���U��y�k���<��>�sK1w�;(�Zp�p�g���w��_�Q�q�a������0�6��S9�.B��L7	2E� )'�^�y�W���Yip���&�Ő�����c*�(�`ԣ#x�6���FuFs�Ro0ȥ�T2]������R���"*A6㯉�\�M�0�� ��Yy��a�M�&h���O���l�&�&�ܺc7�vӻٗu'� �@ը �{�:j�0LXa 3C �<���V0K��k�M�z���ˇ���L�%6`^�C��g*�O�b�hj���t�*6w��d���[�Ӱ*Y�&* �ɇR�h����Ϣ����j���s\:�����m�<�qfvE�L$�RB�a��m�@&�JT���
|�T��
)���E\�7�~=�yD�����!�����)��l\��u�5�p��Y��U��C�)����س��;B���)�|�%p��a�f9���"�q�?�q���*a�c�~��u\EK|����n	��C�*���@�*5�@��K�sL@,����q8x[H�T���in�<PT	��[��hh�|��z��:l#��x!z�^*8͍��Y���e���+IsyY�����(�>7M�VWT��S�CL5���ZoG翬�5u�}4wA԰����,�Y�xt
$�l F��bTwW��53����7"��bc���Hkl��U�q��"
xi$]͓F@��1��!�vQ���wP�B?>`7�H��E�[�6or���p>C.�a�L�<�'·M��:�q@�+����{�k��Oz6�����(�ԛ�暏�
����R���˶�AgG;F���6z]�˂}��f�N�[���_�����v�7)q1�ō�ve��%��Z�ǞtJ/�(��y���@ �^�[������؞m���'��(���ָ6~��[=�Hv�cm�_8���Ҙ�8)�q��w=��t�$��-b�@�����u���y�N���DB�B+�MYE~��,�.ܼ��vnA�\Nnc8x{�� ﻔ�"���8�R-o)+&$WX�Ih�rp�,t��vp@1S���*�����E��S�W�c�kP�DY3�^���+ݟ�ƙ��ז��q��Iْ��8c]��g���?�a�0�f�Ol\�������n
�aU�#�	���|���U�hmzGS���?K�!��A��F�4U-N*'�{/�P���D�z쳞#&`��H�z����pX�4�ڿZ�R`�2�E�m0���\��C�E�1!�s�._�����#Y�~~$P�/ǔ�y���j� |����x*��\/ht���QXh/�α��R��WSRc��Ax<CF��]urn �Ƀ/����k-��m@7%$g5�Z�99b��Rcv����Τ�>|ۜaF�,Ktf"���Ȭ���fq[ ��ː�Z&U������Շć���(�6_�|�"Uw�xp��@����.�Ƨ���6j�z^�[�0��?��xO���Y���'u]�#W�%n�g/x��l�o��y5���}��>0�0�e������qل',M��o��Fr?	~(Jy�7�^M_�y|�4W?���M�Q���Cr�YƖ��8'轨�+զ5�Z�<��͡2����$pw�c�����gI��3��I�8��E�D��� �PP^��������/Vt��W,<k�(G��7,��6��!����A����9��Z-˱<ar��&w��R�����4�W��'�_�/B�.�z�P���IE�9���"ħ�Yp� �ʘ��ߗ�?=��|��;�rI
��? ���\���9;$či�Y�ƃYW	z2Hz��c8�z�K�������&Rٔ��L�>$:il�7Ol���1��!��mն��l�@��we���7�9O��p4e�Vw,Qjq��A����ڍ�Zjy���i�}=S8���ճo���9GHC��n��Q����R�+Z �S:1R1Y����-��jm��S�\��JT�$��a_x�}υ�Yz��
�%���@щ�i�m�u@M�e���S����:�f51k2C�8Q�����m���x`����s�KޡX��ϕ<$Ά��Z:�"���Au�?RV�!���f�%�S�i�X�G7�/Pc�p�a��Q�����d�q�]�c.�g,-�C���ee��԰�
����2�j�U�w�r>5�97�zKd�L���UF�#L3޳K�s£���ĺ�CDa���ű}!�@G7��ӏ#O3���;l���m/S�6�D��o������_U�;ڕbFBׇ|����6�%�-�#��Ta��H9���T��u�ڲN�F��z~{�w�s[��C��|#5����,����%y�4����3�wL���ʼ�;}T_GW�T�{ �}�#~�`��X0}H�#$��K�����͘�h]���T��'�V�,���b��P��6T4�?�����~QN�3����Zwq&��Y�kkO�yg�F�Ճ�^�~SXcRX(�ú"���ݒ����E���\P�Ŷ��bo�>}��Z�WX�0�������c�Xe�N��⪏o���	��O2B�~L�\Z`��2�e@.��Y�؃K[�`e�Vb�Z-�'�|�U�?�l�cfe)����b]�N��I��!�2%(]�!�^*��&�k��ē'�Y�Ԏ�T*�jO�����"$(g� |>.�3�^��Q.��J��A�B��Xp��"��f_���c;"=�T��W'�� �tرZd�є����{
�n�Zs&c��i�OT��@���	�53�P�dO�����W,w��
D���toA�"�f��sx��f6Y3���:d�-��L��k5~9���7uyQ��{��t��z�ө	w�[�����Bh����L��à��͚�Ӟ6^�4��k�HcC�ť��]T1G���%�%X�i�h�z���WX�ֿ*����ԍdΡk]L��`��i���7�-d���q�:|\�:]j�C?���tYhoԕC�
3O�/)�����?��/�G%����{W����&�5=�u��p���N��Y���>?Ⱥ2�8�R�6�ʘTRg�����>{���o��d�1I͌\�,
N�a;$ˑ�R!��I9�,�y &��9�8/]6���c�xq+����>"q��x�F���l}IZ�`�� 5�myQ�M�R 0fU��-�IB�YR�K�g�r8:#��螛�6�r�^�B4ְ��|�/��`���]$nR�R��p����r�ބ��?ɸ�[���cV���E�k�&�%��hJQ����@R��mh?-Z5��1ѣ�K��G�*��.��Em�o~���"])B�{��+����-�@q.�ي�b�9���� ���f�_�G�Z5��Qi^��
{St�'A��vCB���?>
H�@X\�3��;ُ.���YG�A�E�[3m8� q�P�_:��j���?��P�6�=�k�,(���)K"�v��U�T~1(9�%7'M��?�S�U��ދ-`4��EP��'8Ȯ`�eo6���`�D��G^�yL<~*��-���F{��f��x�!^����%����|n�����*n��W�hHGXB	�	�3��xK�AY��[��}�N��n�V��I��,])
�W(��'&�s�1��k�3��'0�[C�������m�:��N_��{��Z'���#&�7ع8T�����i銬��D��ܻ�Eh���@?����9��e$Y4������\�����Y�R��:������
�L�_(z�Ŵ���}�XA|.pS|p(��T9���Z�i���<ޯ�r7o��e/�/�>�)�b\T]ZG�j}8j~�?W"c��Y�l�A��3U�F<����bm.bˀ�{��AOV)���������y���Z�ȭ?�ߜp���ҕ����lY;�/��"��A�x�5�M��k�Uk�n�K�x�B��C����JscQ��p�A�����/Jä��~���Qy�`Ł���SH]^��0�eS����e�!:� �g�L?��`V�.,�N<:^�)�x?�:�����g�������c��Rb������P�z����*�E���k�Th�'������\���=]���25[K��;���Ț7��;��=��s�����Y��}��^���̣�1���b)�����Ӕ�H=�5�b�8�f��1��sN%�\��s{������t���P����[�V�zOn��b���Ȉ_U͗YO���o����,!w(!��.���-�����M���ဨX�Pw�|;*����M�X��'�B?
�5}�����v"+�P��D?o=�S�6���2j{l��~Q_:б�|� �>6�;�1}@�����
Yd�M����\b�Y\x}.m7{>)0.�7�>߰����]z�m��N1���ZK������Y�068j����V}�[e�CT��8�%W,4\�/:�k���~yDDQγ��ln?��Z���G�0TxT�p4b՞���}_ �s��25=�E��D��U "UhO��G�8O^��ٻ������BC�K��[Ƴ����f�S���nѓ��C� m({o�b�8�KnVN�>q�je��H(�#i
�֧��1܊��T�wXB�ʅ_(�&�W1c����8�pl�j~����G�NE��"�V(�} R�vࡰ�f�t��L��whQ��O��
���amP��e;����M',o����@F��Q������>g�-kFU�;<nf����q�,�!���X�e��4��|pY�v��PG:Ýe��c�-ŚUS֨r_�tj0*��^Q\l��?[5R�Z�D���>h���;۱���H�i���_�+2�J����!��ˆ��Mt��_�����>���7��|a��~��wFi�&�j&jL�2�[L9%`!�+�m?.��
4d؏rC� �%��Ҍ�X�SiCb2�\�	3�줨+�zx��r���;�O�;o���"ɱp���A�%%&�~7�4�)2��}��&z��<�-������ܴ 6�5�ְm�Z(7�z�a5��2��'~t'�G �B�c���қ!�a�S���L:�-���ݮΏț���;4�i=+[�>a_����/ Ȓf](���dPm�Y���*f��5-x;����Zm|*tĒ�Ɯ�qٰJ����Ɋ�:<�33���L���0=�V3$�K��T�k9����w�{�o��?0-���f�s;>gD�f��E򂢪�ş9������I� ��FT��v;��G���/�j�s+}Lq�O�>1�)5�<���|;)��	�r��cWB��%}�Y����xl8����(�a��.s�0տ�(5 �@a���Q���| ��͂�'qE�R\G�mj���� k0ۭ�o�J3Hn�mm���-8�p�M��6�hM���EH�^��x�O$��B���m�នN.gę�=|W�^� �sW��;�Z��P���V������i|x-�5���^):RxA	~Ǥ�;ǫ��K��t�&Ԫ�i��`���'�C�̈́�an �,�
�M�+8<r�o�
J<�l�?�(��8�vG��n���wu�؃`�$k��[%�\$�=������u� ��[&l��`�1�Z5ug��\�D&��'2IA�vk`$Y<kPN(�pVb�N	�C�N�Ox��_s+U7}�.Ԋ�5Q�����ז�}#����b��HT*�����@>��p�A���H�pC�&Y~� F"�}U����`��Y�lq��ֺĵ#m�d��)�ar���wQ1n,lOa�{�F,?3��?�l�,�꿬øK��h@ˊw���Н�h?������{DF�R.��$F�ԽtJ��E��x/���r�5m#A�m�k��q�a�.���.P��������$�MaDA�H��I�p�O{{�O�M9����Yjٳy�RЦ�>��`��q{E��k�k����`��'zI�Mt��b�o�q�j�ʀ�'r��T�!�pI�v��o�H��o��x<|��W~9X)��0���@�<CۖR �)�&���P��2+ݚ���Y��
�0,�
��b����O��o�)��V�M�hn5�\��ݧ�s��(I�	厝
��F�V�=�����[���<�� t��S;u�p����S�E���f�`�e�=�w�,^^	��~ы(��B��V�e�I'�?pأ?x��hHZ��f�����p2;�\^��m�������憔*�ek�\��g�XZ���;�7ũ_��=X$ZC��e��U��� �y
�|~͝-Nc'y�7p9�H��"\��Ԗx@	E>咻��Λ��p#�i\,W�_D��?p��d`Cq��P&�������9)�d�3���%W��ܗ�2rMm��|�[��<H���#������mW�nH��c��G� c��d����NEG��DA�5cm�� sC�[R�%��Y�s�d��ϰ��_����%H1M�u�~���i#�`M�ǟ3]7�یڑ�%�>	.�[��'!��̾⨆B�c �$����=n�SA[�PKzZ*T���^������vJ�X*��n��s!"_�0E!�ʇZ^q��n�0����.�-#�D�2D*T��Vzo�����#�|�e��鼙�U����O�!�^���<&(��8����\ߏ'I%�ǆ+d6���Q�v@�b�C���;�X9Z_�7�t�|�L����6.�KM.G���r�BFv/�Q*{���T��o��	��ˁ�̟ȡ��m
2i���-�%co��q'�%����qW���s ~_����9�bk����ו��:u�as�u���v^o[����JPq^�>E;�b#����t*�'m�u(@y������O��"v�|8�Tmī��8L%�s��'��/�X&��r|`v�y���D*h`^���������֊��d27��r�Q�7|������M�I��!O!��%��E���0b�>24�~>������e�1�'�e!��%'��=���=i�R��)!1����s����BRn���fPf��
w��Τu���t��
Q�!�K�)���
�(����?W#��h`�~7�(�.�o<0=)��J�N��"#��fy�� b����õ�g�,k����Gx��."�/{��z�߱ǒ�?�_V�Ê\�St���e�$S�E��!�
�X53��A�3�5�͎��n�흦B�i������x��3ur6?;�VF���� _�,���:P���^�#Z�x{�2�F���JP'�K��dKB��QY���x��I��Xp��k(炠VC��Xh߭���w��g����m���F/K��m�-�%A�kj#4�a��'Xn�����Y*�od�\ē` �>�^9�C��7�1L��[S�V3�<�+E�� 9���,��U�4:f}�����b-q��@h�Wl�"O��}�r+�����{Q#��L�5�Mv*�f���v�NX�@M�k��}���)�����QxcF8��a]:s�V��d_�	G�x�Rp�k�Ã�նt�\�=&h�o��b�I[)/X���^�����.u�)o�+I6�8;Wд���A~��r��Y9Ι~�*�Nl,zԋ5���$��j>��qY&m\�{p��spM(;%3³�\Q9�#� +v���07���cv-C|�>&�jqzNRYi_�9��X�	�̄���.:�ęk�J�DJv	L(,4��� A�{Cp�(�K$-A�',=)�id'a�7��Ìq���<�%�L
c���³���O�#2C�s��D�7[�ϖ[N����SU��c}�E�ȃ�2�ƣ"��<,��Q˧0�J��� ��n�Є5��w��ޜ��g�/N�輨��������4䫙d��j~�u�H䩋^�+|�z��"� �x%p�W��Uၚw������S�_]��L_�٨t'���r������ϑ�A����;�l8����@����� �)JRJ�9��D��2 �l��,�j�� ꭥԵ���G#���q0��M$t��ļ�a[g ����q��z[K.oZ%�_)��mkUG+��H�h�D$��?�<��6�ʨ%�^j�o^��!��+�$�m{u�T�n�+w3�I��Au}:%	jۙ~�4
�@�'�B�:$}ܭՌ-Ye���8��:�w����M_Pc�r���c�'#+3-�	<<�y,��B��b� 8t���tz�e0}6%���'y��J��6�-�wH!�|4���3M�@����T�鎚���Y�� �~���z��_�d�1��ʟ��`q���XH;��YbNG���8/���:!v�����Q��>�!�"�'`�r6��s���mH��Ӧ��7M��?Ѧ����":��>����V�k�g�M���~|LlL�o{�Fjk���Т���4%�zYB�����f�wH�w�q4��O�C5�U3��k���[nw2����V���������٪�S�����mZE��؃~�JAy'��8Tӊq��r�M�/���L�hn�e�O ��<EѤ�ݬ�-kd�*M*�&�VƯ��m�(jfI����1s�������r�d�@�{�Hx>!ؖX���k��*�a�80R�l� �� ��@2��4�T�{��!m8�)��<+ꤪǥ��qWs%3WX��;���L�CG}��I?����qU�Z��u���ΰD��Y��{������H��P�D����2��}��6�WN��"JY��(����j���C�ǧM�W���QfT�=V4�z�[�xH��A�9,�� ����q���%x<�� ��j�#D��g���dޭJ�R���rܓ��[+�f�&�z�8����������k|�T���eH��)�6j���*������"��E-��l�=�D!������\@+��4��B��|P;g
C��Y���\.X��^/��8Լ���W�R9^��Ζ��~d�l��gp�����**ۀ���bQۉ�`�C�' ��5-�j��N���d�vݔ�/��jgd���6쀃��0�UAk�2�6���)�_��&���,ǉM28͗AC}�������Zpw>`�}~�U�0��x��y�P6������H/�f�D�~���Wg`$$����I��Bi��lj^K �Ҝ����u�{�'p����*�E��7�4�UmA��Eh@��qy���
��M��~��}Q�
��}w@B�H�C+�@=��k8L�IR6W9�|����N�}t�[���}��Y�ɄZ�:S�= _5����qa�Kb`,J�^�H��l��4�\W�Sg�'��cq�uIg����@(��ɳn=	�_�e��v��P�ٛ�'Mr�V(oHO!����rb�[5��S���LpZ�Aۜ�%WhB0ʛ�r��>� ʺ�������ye�ѹ����������W��^�4��4�|ו�ڗ�;ԁp��>�9ke�,!{\�7�!M��Vr�}q�,rI��WN�k)䗛B6�>�`��0�n|&�cYP_%㯣v�,��$E1�q�,œ�Ք,����T���B���v��A�>�$й��qC���yORʴ��.�����P����}�CH��w$��y��`ى6ts�Nl����S���� ��9��K䏖�F%:g��1�z�)mz������H%�y ��c,]8�5��y�Bp����z�۱s�f=�o(��	b~3>��8	֔��Y�K�C;2=P��Y�^���c �3�MX�[Ϥ�ݙ�GN��.� ՠ�����LC�����Z�U�0d�z�0??���8��Im��C�F*����4�Bѹ�̿16) K���qJ��Z�L���loY�$C�}�?%��X�hU�e
��E
�Q߂v62�tDd8㽱�8�yj�7��� ����$:, A�m��f�\{4ôJ��x-S1�3X i� ��6P�N�:���`-q~T&M��"+3�����;s�G�}SX* Ɗ�+��Ꮞ�}Z�VKdE���gTJ)*�y�оw��@�=��<�i( j���.)o?��֡ H�W��b���꜖"ڥ��G��3�t���=C�W��v:Y9!��eݲ��K���==XuǸ�1H^���!,KG1�����x"8C�6OY�a=k'����o�n���8��{�*n�q-cܗ�2�8⸜� �I�h T�W��=�����LR���b�تa�f���nt�G�I��~ꝧ9�j�e�-\�O\/h��9��鴄єPj��kFy�RH{�$IOX������&v��Aƪ#:�x�p���x�Yx֏#-Zy�����$���v;1gbC�z����Рg��������P�+D�7��$���{!Τ�V(R�`�ܪ2���y��W����G���I���u�'_�rIb�-V<��Iî�X�-�4e|3e�O��j���<��pa6��=���h�,Y�ic�#X����f�����&��v����{={O������I�%
e��\�z�67�I���m��ϳ=���:���<��N& �䯌=ك���.�߮�i�ii��TbD�"l�q�'BS�6��,.
��u���mT��������~7��0�sn�K�2?�hs�������typy�
�%��!�5����#>�;ܩ��hE'�#6���K�H!HpE������
�C&~,��HA�Y'y>�&n1�� SAW�`�o�S듋Ps��q_ ���#��́D,�I���-����?�X�2+��Z�3�q`iF�R���5��_�ǭ�.�.�X�u���8�[]�f��z�9���儛� �
�Q��v�3��k��I�����0�N^�/��|��G�T��C�!��%�6�-�$������G�Zʳ������q�š,�����9\Uk
�"E�&���o��h����;Aw.�c���o��t?�?mMtu��r��,�gÒf[�9�ͳH��N_z�nL��W��E<NRU*G���#�SL���1��~��O�v�#���)�@�%�r*e��Q�2�����L�,u�Q�+� T���¢fF�E$�DbȜ���9l��+A	Yn��I���~\���.�����Y�C��/&��Gn�~��n=�h�lNkM��s�-�E�&q[?.�3�Ek��`}�Q����ӈs�n�ዛ�賅u��8�N/u��ڗ�����&a��s�U���,��Ǭ;"����J�����#���C2�9�,� �����YM;kl��/�'�B7�ɢKː;�q�� B�Oq3Y�U}��H���g��!�'x��ޑ�O�T�zl:�,��.F���rd\�0|3�;�&�ߪ�KT�Rm~:��j,�� ΐ{$hLj�͵E�[��j!����.+B��?� ��C=�?�lХ��N��KRq�uϷi�曁�J��J�l��+��O��LԳT��W /Qd.���}����M[�â�ҫC��)�s��,��A���)ԼR��>��r��ָѿ���TNM���\���gB��4.�OYb�j@O�n��x��8+����1�h_�|`�d!2����"¾�kI�\�8���o*�d\�B�K"�~�φ��K���|��g�э��d�Q��D�d���W��I�!�c����O�_;�'�ш�9JQR
mR����@���ةR�h�Jy�����p���vW���[6�0g�)̫%��/�U�µ��0D�a��T#��u)l��)5���0���������e��b�����^�Y���
�V&�戗)n^�kV�T/��Mz۲+kt��3�lr��`fx���/���Z�m�>5"Ru`�;BUG�5r�8��F�$� ����s�>;P3���!�=���uL��������E�	�@�o���y��:2��T;K���]]g-�3J:�{�D�|a��1x�&�8�Ԍcq�G��ւ�<��� .:AG	�R���v��v�P�Ȝ��F4�K�` \X� ������co.H-�x���~���S��}8$/7lw`��"����<	/�@�;8����X©������q����C,��ؓ2a��(]��w�Ҙ�W�I�@�A�4FD��0Uo,��[R��Z=���7��m�,A6�F��D*�47%͐28���I~��{�I�E)��֨K/e�-��Ӝ�{L��]�Nڽ��OԞ1�{�:L#����z����Nc��}���6�$�)��%�rr@ڙ	B������#��Jm)s��z��%-SK(�K",Ϋ���X�Ad65���2�H|r9�4-dx�s.dcʾ�Ь5'ѓc�)&@�K��m8 ����L�c�v]��
�v�[o-�eA�
�")`ݔ��<�I6��AkN�<��t���	�\P��&m���2�P�w�=����蒷���IY�����f[�HͲ�HS�e%��v��}���~G�p-����GǬIi-<%�y��	)y�wJH�!䱭�!{�,�.��@���D����3H��;�2?�I�0Ո�����gf׺7s@�t�eѫ�&Լ�<��u�J%gґ
��S77���լ��k":�O��r�jiDf'���T�}���#���� x���J� =��)�q�#�SM�a�D0I_��))���o�utPul��L:"�"@���} �!�UPeŭ�3��Q
���Դ{�)1\>A��˦2;��ݣ7��^�!c�P�o��0�'�M�;#_�"�>k���:�T�?RJ�p���*0���ej�Ⓡ� 
D�bQVkS�Y����%~�'p nr^(��̐��F
��8J��>3/���q���š�*�%��N���6yQv��w�>#�:k{'�`���`�l�ܽ5�V���7a
��k��;�~#%z:q����h���G2�}Kn�r��Tڋ~rw��O0�t�4��+F�)i3�i�ͣ-��,��ʭd��j��|����%�x��2d��ً�֒�H_���І^�
s4���Z[�g�v����eA�u�{{�S�Q:>8����0��.p��Ϸ[L�E�C0{Y�]��6A%]X��8�'|�ė���k^YS�4�ZZ��W�mwk�SRcs4ۣ�[�i�W	8��5�gG�lH<��d��g�C���B���ϕ����0K�1q�&*�}͌��fg��Y���&!��4�m�B!�S�ɒ�訠ޞ>R,�5fHʜ^��#���hQ<� b5�A�ց�U��3�H�բ8-˒b��^���t�4��2���K:�O��hѢ_�����C��!s�l���{@rM�'��7eH��`�<w��`�2Vd|���zϪ�^��W]Lx[�4z캕�g�+r��t��}\K�kHI|�w���MԺ%4�y�-΋o�Ye���#�����"5�4��*�����"��K��G�?��c�.o�Js1HB�G����b�
�GZ�o[�J��JT���>3��z&��A�ڷ�K��U������FW93i�W.&�91����-�Q�<'����F�ه���/�rdB1���p���"���'nzr���),Ŝt����b��M�i�#Ά<9�{�~�R���9���(��O�t��JD�6�Z�l���:�ؓ���giĽON�}���[�T���&S>M��N*����1�:5}QT��:�{pʺ��A57ۧ�n3�W��mh�����1Mo`3��]#� L�������-:=���l �y�k�ͱ�=�vo�U�w��!e���p��Ѹ>������w�RK��]���gt3�l���1m,�꼑�;)�?�,�\�Z2�����8�6&O{+E�ȉ�B0�?T3�i3HU@�XE���7~U����_�XH�c dǛf4��owr�k��h�L�l�C�j��tLn9��z���͔�=��˿{"+����M�-C�c|e-Vo���vŠ�|�Du�X����|*Rʜ)Ihl3�X5*z̄Q��n��l�QZ_���¹���a�-2B�i��$G5�2�p�������5��ip��U�d,���b�� f��2.plo�U>F����:Y
]��
l0��l�(�Mb��8��̴Cb�0�;oݽ��tX�L�G{]	f�_	h�jP�$M�|.?��_����?�2t�ˋ�>�3���"5��Z�&k�EV N�4��������$bzTxؤ�������R��'�^����iO��t��k[4�r��Ķ�-�TX���K��m��6b^e�d%B���ܒZұ����t��7�����"C�s�_	�&��7A�t��=����z��{�f ;5[	�ͭ�!*n��ϥ>P��|}A�H�3(����L��3��|��d��Z��׭v�y�������hl�B��F�YZ���(ީ3��;��~�T�z�[�H!JHCO-"I�- {���.)/vW6���z���Q��m���j��mC1�=�ò9�8<{Wɸ��Zs��/�ɣ�>T|?o5��<w����@�(qƷ���"S�j���܆�i�k_�l柉�L�0� ���g�]<h|�����׏�L��r��Dߘ["E(;$l�w�l��^�(�F�emc��\5b������-P&7�|ě�t��>x(+�ݸ�Leь��,����h�kCQ����$�%��	r�<�\�oX���*�p��h��l���Eq�����l�������u �u�p�RI��K<�����>�gv�H��8kc�/��
���TYe���+�F�GDs:{q�wܴ�?�V��->�������uL�C4<�!��Y�E��84����U���0Z�hd����Ai����{0	F�R%a �B�ʜ��f4���\c���?>cb�>4�7Hy99>,�OG�3�	+G�A��^�I�b�>�&O.�&�����|�.bW��r���{��4����yd�> ��<�J�,��,��c߭����5S�A%�Q����n�
m�<���]�^�Xt����~��X�K..(߅���F|�0�͟�g܍�<.T�Z��\$1�2�诹�� C٤���٩�t��n������I��p��җ�/ rЛ�v����a4սY��X���c���}�Z#�d�8����E���v_�f|��+f��0����	x�R_�8s��lF�C�z��_٬�V�fu�X���bʦ/�<Ɵ�]���(��+Y$��Zh0O����:�h�b��[����|�'q�A�*��ב��"�*��~��Y�����I^g�����^�0� ��a߷��Җ=��dX��I�E/���M���r��G�ma������¥I\��kN�o�qA4L�;W��h��8}�/����P.-��+/���_& ��G�x�ZR.��++��ߊ����e<�,�l£��!�䩫���C�7�]����A-��K"�
�|�1���n"xNW$[�6j�,�ǻ*}�����֔�3bu����"��@="IU}�����tDW������7���B���0��x?ϵ"�D�~љi�(1'GxF�(؆��@E^����GJ7;.�w?0�z���ZR/���z����s/#�R���HeA��^��G�kk����R挭s~*���ln���^x�6�#���1�N�~�c)l���o��Jrvl�0��%~j�ۙ�KXƳ��܃������ϙ�H�ɦ�~�g�Q���4�72B�ޭ�C�<t���>��gH�d��M٘į�Ƃĺ�0�$��l"�,�V?�ٹ�2jW��#��~����!m���m�����c�P9��w;l�]�������;�pF9��|S96=8|A�r@��M �׋���cm?$E0���_�#�� R�QW��-�-�3��9�	&�/�o�0������)��C�f�uÓP�(��S����c�!��v;�s��sŃGp��V(M
�q�T:�����4'���*��ҏ!܁Ƥ&E�8V��4}`�|<�9�t�l�������/�&�L�U�$+`Pi�|����n�w%'
��I�J��1���O��Cw{ ����F3j����dA}�.�f1�*Wp2*�El�p�z�@�UO�K�W�'}I����/k~ڟ��V���v�����a{vaῧe�k9Q��~k�ۖ˵�v�[���u�9�-�N�>rT���h�?��W��DQ7ԅ����Q�������Q�/�Qe�6��)�U�ޗ�3��[�3ԝ���W;`N�,�K��g.K�6�W��t��^�R��̪q��t|�K������:\���x�Q!s0���OB�tu�cO�.'��x�T��&(� �R�^pۂ��`����xz�g�y�����E�C&�C��L���˥�O���4����ߒ{�/�-J����.����������i�
�7`���fj�m�7G ��x�YD�'y��y&М��;�O8�ʇ����%Ss��0�W����6$�p}��/hH�s=cS�v��f����0iZ-W:Α�P�V�xg�e�zz��ɚ��R��Z��}��9�G4���	���	�`�>�A���W��ٓ���ɝ�Ѷq���Y����%����k�%��閻�v,X&��0n��en\���ʶZ��1*p�g�%҂�-|�e���}ܴ��Yt�!�&��x:'SEZ�x ]�ي���Ó��5��l~��F���UrHJV���^a�Y�9��*ٟ��	�R�`�:���W�����!�?�|���G� ;�82����"E���^�!�u�t޼�cV����e� ��	��hc�2�3��'z�akU�>#�X�iQ�@u	9l;�U�~p�5�8ek1��	�c�#�	����������'�p;�ۣz��a�m�Aф}����<��>���@�kwm�{��\�ƶ�$�q�n#����~�UI�{�B������.<kLf�;ZO�2#zK��j��=��N�{�8˒�i9S�.3��1xK7_��6�i����6�5��=�SAGG�����v��K��L@&�|��MKiv�	�
avB>���g]6��,���c5�@&?�����x��9��ط�f��+ ��3�p�+2�Bm��	O2���� u�m�	��f�"�NP�Yv�"�\�œ�41j��L���l�6C�S�a� ۍ�))PwO	l��hJڀ�;�`����y��ax+��&�.������Bݜ����+�u�L����K�w�W���-L�g_-Ȍsa���P�V/bKX@�\�ΣB�Z���s���C��:�4���ma���y?YԹ������̀ٗM�S��Ʒ9,�T��� ��h�$���n�����F&!�e=�3�~@Č��-��8�nd@�,���U�b�t1r�z� �i�vM��1�	��6fj�;�@=m!Ҵ)����=�*��	]MG#�i���^jJ�0c
X}G�X$�P_'(��V�/������ٕ�ۺ��-*9�s�ԁ�=�F��L.O�߻�b+��2���������Kx��*�|	��\[}yxY1����"���jfR8[���E�ߘT8�]��[�l�u®#���A�Zp
�B��-�kLB:��呎�H��u3�Y��3���w���A�$��*����qpg԰���=ǈ[a!�Q4�U����{����dI�q9d��Z��ς��J�i!{,<a��`�����3�ș�9I�dI�`�<o�H/�K9vg|���QWgD[-G_�����V����}N����ӊ���ʠFe~���Ց�\s�5e�krE��N��E6�k��b�`	��gNx��SPk�����Ԯj�������^h��G�����+y��tU#��ز�u���� ��Քb�tg������t�\mD�"Є�C�@1��X�vn ���-"�潔�?�A�2&Յ�*��Dx���YD�\9���f�5?���cA�w*����f�+_?~����M10s\ &�S@l�+5�A�L�Px�'1���P�ڞ�f\��W��=N�j���&(UFf -�����}�w}3��qn5d�,������c�Xc:6qO���z�*OKS��E]o4����_Ͱ�s+d+��)��k��
�F��h6I�Rpk�8l���j�6QOf!�L�
�;��_n6�����`����,S d�H�A{i�0a+@��/�SRW�i�������
@|P��N�p�7��ݜ%�H�:�oK���{wE�1�^��'U�m�a4�M��f������-�>(~\�����>���\?g�i;��cռw%�_Y�*r������Qe�֩S�-*9��b�[<�0G��b��g�F�|��zt"68)�~�䟟,���Ũ~a�s�� pt�0ʞv�2���d������w��_!��@�>�LC%��yev��Bϔ�EY>.� �sY�֥Gہ�r{�bʾ���	����㥩Ҷ'���濋c�� ���,D��F��5�?<��Aҙ��[x��V*���ǎ`>R�Ҥ���� M�<�h�R�aӤE8�+c~o��uظ��US�N��6m}A@'d ��Y�lt��C�E	�Nߥ�y��*`Lxn��}��k9��ܔF�4�ј����E ��`����@�V�M��FR�F�"�U���Ȳ�ޱ��K	��"A��	FDH����c���'�@�Mn��[&$��F,W�OF��ڱ�7dw!*E8̕�K�8�0���W@\��<�<)yn��w�nx7�v�[ƛ����y��c/ť�"���<���x�s�,�M���r���˯A�&���Nђ��|蒃�ov����Ud?���B�9J2S��&<������C1�,��Q���^�M�w������h�@pmR�>������A�x�� ѥ~����">K�G<��V����g
�Բ�3�_ ��lD�֊X�ez}f�S��NW�O��y�e����V�#�=%�y=
�s3!ۢ~�P2R�� 1�M�_�2F߁�3�Xo	;W�;�o���Ju?��3����G&��"_�$�fYd��S�H�vK��a�Vm{���ŕ����A����gw�v�ǿ��1� �"V�E7�9zǺ x�]M/7����~�z%h��)}}~���U���Ow���#��p����<��?� }�J%��Y�;�ͅ�N�V�h2/�W��
�z��e"J��pz�~��(0�w���#�R��م�l���ІW�SB	���K\��qS�O�/_���W�1	���:U��W�o����H��=c��ڊ?��?����e#�0ol��5�eW�L�;yv�3�7d��ocT�g����a���"�6
�[/�����S9�;5c���9,��-�&���~�۽��R���Yi;�h���XI��Pj)^�\��}���4f�c2Q����	�����׺�*	^$Sk��:��A �ڣ�9�2]�6h���Q���s ���b����`��,�u5_N��D��,����=áԂM��-��a����RXX{?�wo�^�)D�%����h֞3�N�������8�R"R�8~X����Z�9�-+�;���A�x���я,������D]�DdH>��QM�au���(!_�GVin#�qav�82������"ȴs[�aOg\^�[��N�d�����#Kxo�Q�J����"�x~ �����q�)��Q��eq�I'�,ި%��Tva���3+قl��/�1�W�P�].՚xG���_15�� �yn���3��(Er���W�s�)K3KU��O��Q>O~T6�)2XQ���0*�\�wZiTn�霿g��9��m�*n%�Y�����t�m�-ӟY�i���Є����k?{�"�T�^��sTd�Q�j��$�b���5Ä#��c2����W;�.Z�`�{͍nnߣ� �#B6��sJ�XC�6\�`���G�Q�v�J�^�ɲ�Zs�m�eýL�Op�B[�,��3j�� �q�0��}��?.�o��|�th'�;a)�nn�ۓ�WU9�-{�ĥ����Q���'\��&�:Ri��ms��Vi[���p�I�֩��9��� �v������9_6�]Q��P�u��9�����X��擙,�F�e�?��6�Ӵ���83yp���H�EH��S`L!�%SM<F�:�ꄷ\��W��96"�/�
�����@�^�m[6�A�c`h����LI���dJ�jQƬ���8ނ�gP1��.-C�����7-_���ȿ�!F����$��J�����dT�8���6GMp���[�*q
����9�T"oW���%#I=G���
���B�Lt� ��g�'��q���A�	�cb�ٰ �屔�ő�'������=ƫ�U�i��<���꽲L%}�����8*"�������B��ߗ�1�m�9��֕�g���)��yѱ�\����~�:��^�i���2��0���#j�ɤ�>knday2��qK�=*����	b;�y�+�w�%��<�<�Y�[\b8��L��̄���ODb���� Ә�:_�X��}�6�xʪgM��.��g*���2b��劖1+����≢�$���:)E�������h���-�(��XA���ҙ?(�D��`#(~��d�����\���X�|��O�"�%J�#Nh���A*Wʄ��b��F�-p>!`b��,�Ƙ�B*�k�J2����a��1���� �c��Q�dþ_δE�piZU4�˅>f���aԴ>���2�îٮ'H�)߁?��7�DM�1Ķ$��jN���$b�H�����B�0XfG���H�/%k�7�\2,�>|�8I����F�����$$g��� ���c.D���`s��(( k�#���ll����l��ci9��d���'nd�˔g�Հ��!Hp A-�E��k��8tZ `Ց��j��M��3��}{f���$�9��Ye�τ^���oߴ�/������"� ���V��$�3.�AHl�.q����N����$b���`� ��L9�����>{�	��렊��3W�!.u�"�S��4^������W�O+���b��)���:��."�����	��d=X\���DfA�,ԠYb d�Ԛ���+��_3S�O���9F��94ett�c��c/�ŝ�i �!C��j��A��-�b���ur�j�vA�Kq�h�����Se�1�hV�Q7>�"�l�nuR���2	�h�*��Ĥ>�j�II+�6�Q�'�KpX`BqJ��U��i��y���+� +>-`�A��Α�IMn�]�k��p>,/Ѣɍ#�
�έv�sqR?���E4S�oZ	�Qg��mW��)$��𸚝�+��` ��ɷb�Е�	�&N����0���fQ�w�u 
�f11Iy�me�,�t��j�{:S�o�a�X�k�h9�#���Y�Y�F*K�,�����n�R|�kH�ȧ�uBZ3�>N�a��O������B������v��ʺ�/^<�9�ɾYIF����P��68���x؝��}�Q,���t��tZP>���؛�e���w$j�N�Xca�oGl�+��Ͽ<����(�j�J�E?����m�W\JdK�K/m͑s���𡎎��~���^��B�
��DhBO�\Jgϳ;2���6��7�(��T��x;��)mI2�2��&�0��s�s$,�:�V�ʝ%ѣZ��k_C���J�OV�L����Wd#Z/}:Wr�<
\D�N��c�M���Fm�%���T�����=�ZG�G�àI��W_9� 9�Z�s��� Fɸ�ۆ�"jz�/�xQ��t�?��q$^�&��a�T�g�G��o�F�Ax@s�0f�䞐�0�"F}�G���I��3�c�D�/[n1暙�(�+տ���3�jP�O��8����>�<G!7a#vs��]#��{�2$���T��S0���y��C�qf[�����?��C���B����(�fĈ�_-�Y.�/���MK?�ˢ�w��F�nV�5��Wd)X@Nf���F'd�x�Ƚ�L������3"���'���M��z|����S ��5�	�1�6:���2k戯��	}��ZϦ��3�v�f�d|M���ɕբ�(��o����h�-��W� �wEOD7ͮ������D��	���!����4��_'��R��{i�/FQll1�(�dX�� 
фLr ���3� -)�#z�Y����.ס��q���1���ߚ�s����	�Z�l��=�	�`�:�"��;_�U�R�����W��3�e�c�����ǮζpE�DQ7��d�?S9\@�;������Ҏ�Y�[����W�)�p����FSV�K=�[�5����=oF[�׍d�D�>�S�G�4~��[+n1��/���0�,D����)O�U[��",��6T�ݾ�Y�@ 4ab~�����2�4��<��BE�\���:Ux>��8y<�从a�T�+�o�&&L5�0��a�:��Bx�-�V�����M� ���X��g�RwW��R��^�K�sh*StϢ78 �r�_����)$"�dژ������(�͔��@� u�n�R(���0՛|����Ϣ-�J���C�5�~ȸ@�Í�H
���gd3
J�/?�����c�o[֦��(hEb#�qVY����ߓ�1XF)AC�g���Q
CWeW-�_�1P��+�Žc]��L�m��m�-;B�y�*k��ڧ�\�e3��k���zPv��ҍNE�ʥ�ܴH���N�B1)Wķ�� ��_�cg!��Z���4���v	0�<�Lx���3�>*	��ý�c���->Q���e+,|9W@��fI)A"�Q��	Jڋm;�h�!{zR{����f�{a1f�~ö�+߹ŷ"���%������Bz�I�8%>2�m�<��Pk�l�w8}��w-�X�O��9�w�h[J�%뙩�9�pLo�{?�Ó0�����y�j4#� ��gK7���pt7��J�҇ft�u�c�9��D�T�IF5�TLz�hb�n"j�Vv�\4f���X�Dd��ba��X�Sn��W{<z�ځ�N@�����a#��qm�ƅ �-�J�U	Qu3D"`^j_P?���;b�D�S0�cNHլ��%���s0Y����!0B:�J" a� �����4=ʝ��5밟vQ8BK�Oik݃WͶݵ��1�7��!K#�SFg��q��;[��[��Ɩ�eh�����3I����@ִ����m�u8\�T�~yJ6S\���$~I1>p��*A��ZN�d�m��M*e��V�ʖu���0���So�g��0��"`��%VD�pO�idT���'&x,�Y�i0߆�ꢣbu�}V�z�-�]બ���X`���ꁥ�e��#�Ip�{�g0L܏&���%��Xp�G��S�`Q��oBc�ev�g�eW2���y^T�Q�oo���Y]����O�@G���X,\�Ab3Z��бդ�C��`�An���!Y�6&�Nj���}����1�s�#I��-��8T&R2ۜnU�:爄��5�|Y\��l��<d}�c�йO�wg �¨[U���� ������� �#=�Y�*(������6م�]��NF���d��)L��`�k�ݪ��\�������;���!�e�*H�����#�f�1�
6�q�A�_Z9�X�T�qy��/�EV����f�%(F��#��+�"d�x
h�~��Qi3�l ��?\1	 ���^�~�f�<ߦ��-��0�Yr���g]��5� �Ҏ��u�����#�K��&�VKi5T=��o��Y~*�sH�2�*<ZA�h�	���k�Y�[��覤�*M���z*a���eΤ���$���Q�ߜ���:��$����	2̊�H�t'�|��<FxK �|���A{����n�6�|הk:�N�(A����ހ�JX��8�YN�J�L������8����v8���Kv\�`�H�FVX�2�Bq�5�T�,b����h��a]��f.�Z��>�JR����?����/����d�N�+?Vd1Ĳ��� ����ߠ�T�!d���C��9.�>ح�!{��H@f�*�t�N�G�0�4xwJ#�~M�Z���Q�ǡ��A1�͟N-{�5ބ~t�0XX�|i����+��f��@�܉��v�pw{Z�눝!�) � P�f��M�m�/�|}܃O���,QF:*��#9JQ����j��K�y�ӊ�L�u�L=������L�V�5:��/�4�wj�;Q0��k�T��>2�X/�ܪ��@c=h�~Kv��cU�J�9�)>��԰�u�+3���82N4NuA{���H�B#��ǝy�WQ���|�N\}!��L/61�����@ҙ�3�|�&�nh�	����^-��C�d`/�˭L�L����:h��A�n�����1��G寑4���q�٣��X�L��Z�M��솏 d%kz� �t4~��J"���k��7�O��>��x-�%>�,���!z}v
�ʨ�b�#��lh|[�������6?�ץK��t�6'�t�����<��d���:��e�ϖ��'8�!�n���)�w]��mr^���O6E��-���dI��7a��.Ew�T�2��m�5qvh�~!j�;@��I	�.'�)�y�K��6Aά����`C�5������\�n9`�|��D1�V�$��z�=sQBTB����X�_s�f=6�*O�z7�8�g��&�EZYY��k{g=�FP�f�E�NQ���3�/�W�ρ�Kv7��AK�X跮�����������-��6#���o�K� ތ8m����cn�o�a�|���2\��ѻ;\�{��fK�e���$��A�s�ԕ��}���k埉������v^����u�̖o1�w5�.� �r!�:����&��$�Wx3�1R
Ws��h#������Sh�уKa0�N�(�%;%�݌0`��Oڪ�QLfl�rR-��#�%pݜ��'흪	Ro����an��f�L�H�|Y��
� H�,�Zyϝ�v%S�3�J�7n�X�F�zJ��#�t����X������\��}d�Pq�'Dw���Y�����K�LOJ@20��~�G
����?�^�ʏVM)$�A���4TBxz׻WF�y�E
T��_���o�w@ĵ�Q�>Z��X%��D؅����,*VN4'+A�����k�����P��1�"i�3�}�@�\ű7�n7��%$�;r�p�#�iʪa�Tb�2W�5P6R[��{�A��VR�kG*�=.q�l\�~��D`���ϴѷ�`�u,'y���8��bs ZݠyS��B1-z���̇<���!�$�w��m�6�o��t�J����J!�"-y}�cCa�Bb_�i���P���)b*G��w�$6�*<t�y�7mJEЈu�@T@$�Wq�Hqb��O#}� U�D;e2��YLn`�Ao�%�S`1�� � ��Z��c�&��zy�!�%o�钸%8`������*@X9��8Xַ�D��O����`L
D[ٱ�$�!Ճ~�Ժ[��~?�YH������(PPZ�c~��U���S�l̋|n�7o��%g��xa��O��F����M�D�쓆35������u�I����s.�]���T7}�R��*Ji��?��e�̾��'���#)����#���֚���>�9o� �e�~��t�P��H,M��e�}b<�0�����*�¾�>ۇ+�f��d�2��B�c��Ԇ����(nWC��3�tﷱW���>19�\q!Tc�$r8hAX.��*�aQ�1��ƫ�E{��U(��f����$[��bA�(V���O�C`'��l�(�0���^Ϫ��~w<��T>�LV��~���������dA��/����za���K��;���y��v�*;n.<���Q�x�U(ś����G�T�:Y�>sX����5�P��i�eA
�B�.��P�u�I�3玻w�kP���#���CE�ڝ��;)c��P@��Z[�x�V%L��|��''=��v �ra�}eq����j֣�b�ZFA�S�t�4-W���>��x��#�������K0~�A�l��D��uG}�Q1�����E�;[u���_�˽�lh�)����}��U@���#G��%�C�N�P�a�ˌ*ߐ}��t��!����I���4]�OsḮ�g@I[�ڿ]}���Q�1J]��^G������r���ꦛ�(}񻳆軿���zX� ����۳���J���I��.�)���/���+x��U(�ŗ롺%K�-���Z��5|9��Lµ��aǭ߭�#B�د��3bhb4���[VS�~v�f�|��9�"t�V]3W&1�-��d�}�Y[��o�5�M!��|{9�����ɚ.<T1�[C˥#p˯xX�M$?��̨.�s� �}29Fs�tG��� J�5��[�z�V�1ወ+N�9����#m��9��,�?���aO�����s��1�~�zB�M���5yQ׳
ԹH����f� @xđ��[j�;����9	���FaY��rI�Z?��V���K�mD�Lb��R��uX� �X�9u����3M/j����NKm��ʃyO�EÊ��_r�F�g���>o����<u��IK���7�9 �5�nQ��!Az���M)��v�R:9!��
\��%1؞� ����ΐ�Wbw#\B�*L1�h^�&sm8O4h��$����������X'�y�-�����.�j?&�Q-��o�}�dnĔ��v> �%<�&�LE��oݷsY�* 8���^�k�N�d##�qH�W������N��)&g}�4I�7md��*�Y�j�3_��$���!�D�Uw��s��z�;��X�<�׾c��ZKm���AHjm�'����B�L��� �����ő�Qs5��������ү��#���~˩Ľ�b�����/ zq�ȑ���W��7v�'8˗��;�y+U��EH$�B�w�OUg K6��5F�%'���1t<�'�t�@�����i���>��,4�����d*r'�G0��%��B����GTB��T3Kq\.i�L.�D�B�>^�{�6*A�M�vD�F�����L�[��i&��ӆ&�"����._n�H/�ͣ� H�c6
������`F�ûb�����Il���!e�����p�V+h�=�x�� ]��h`� �N����>#�T��>�.�����T���gB�}���gL�Y�"YP���i!eIs��vn)L���q�=���aD~k��Cj�}:�@Ř!�3���-d�HP��'�u��g����$���όꃃ�5b��9'�V��{dR�RZ�LG#�c�[lT���x!�go 1�]��������13�$<Q�V"�h<�X��k l{18��{�P��*"����g���Ӂ�[�,�"��$�{��~_ٲ������&ɘ�-~!���"Y����S���