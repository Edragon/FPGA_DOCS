��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`nE`{`��u*���:�P� � ��ċ�vq��� 3������V�MY��mkN�n!�%@^��|�0���U	#�V�j*P�e$����wA
��M�#����`݇8�&��V#��A�Ct=��@A��_��;L����[V+�F*g�zr������cQ�U��`t�~���~��Yz��G�r*0W."0�_���o�`����ԪEQ�9��jH�H��ȝ�t����k�]��R�EL� G�>~*iV��ڵO�(
\�S�V�T�4�Lv(���[��5�ƠC%%�k.+�n�� ���j{�|v�W���D��Y!�����gn���j֦�(��r������W����vׅ�P�m�sA���]�G?h�|�+J��6-I���[��|ޓx��߽:"�  �� �H��2�zs5�ʟ$qŪ<R�0�H��"�u���Mՙ߬@C���S�E� �ڈ�𬤹1TE�FT����������w*65����+���C�ԧ"Ui�R>� Wnˉ����9�h���Z�oZԚ�X��_Cv\O�1O\*U���0��ە�f���f��3�P�vӃ�Q��+#q��Q<��i����}��^{�њ�ER�%j*��rIx
J��y=�ME�W�ع���b^�"�`7�1�'q�ڝ�p�h�Po��T���_[���F�rp�%{��0j����h'J�ZeSo*�=���;�1�y3�Jt��$0�S�?��:@��ĭU;�n#�n�1S�}[��ꮾ{���	����l�C�晡##�<�$������s�b��D�D� , �Dk)��3�%lHD0�]<z� �G�@?_l����Ť�M��,��nR�j##��G����j �q>P�0��۸�����]�.+"�=�����7�e���Y����%�����giѕ��4�'���l�9��?G���='��H9v�j��I@�G!�Sq��Ѐ� Mn [;�� }4�g���v9t�%QY�8s��E����z��}�{c����))�_�LP��w	^��Lvë��y����m�n��%Qd]���y����ె_�v�O�.2C�.)*���*+
��Y4iY��3CϞz�K4�ץ��M{���i6wؼa)Q�EP��Q޸�#Q���E�]]}s�\�u�A��̶�^[ K���J�"���z��Gp�:�`�"�9����?dM!prm"��m�]I�P����u�Kt��5���g�̯Dz�7kAf��@�aa*�Z׽G�yOV\˯Ŋ�p�MsX9�K7�م{�8����z��1 {�(�x���w�Ӏ|7����c��?�ǹ��$���oɵ0W`�I����6�i�����5����pU�	"�AlL���7�M����K`K��F���k�Ef|a7qu�Y�d%���[)��+�_�#S��7�[�A���dL�zd	A+�<|7ה��3��D3�;��6Hsڽ���c)�A�m,��S�m3l�H7xwi�C۪��:an��I �ʧ�d�R����v�q��h�Se�(����ъ�qkKoi� đ�l�|ּ�ܪ$��%��]�╧J�� ��m�<n��-���d���kU�,^O�8�)�`��a�n	Kv��X2�w�$����w^rk�re��M؃�+��&=��>zUp�� C5�IM��E{��r��2��&$��I0&�|;�,W/�q�~�p���� �6���/����jQ@�|�]R^Öp���{)�<
U��7V\�)�����U�.��pՀ����O��^�O\���fc�I}������(V�RaٷT*l���(;	�Yw�Ɵ�b��������ͽ6+���
��Q���v]�	R2){�yG�D׼[�]b�1�C0XQ��7H� ��g�� �k>���K.��<om`G��|� A@��f4�ԩ-��qCt^[�I�V�M�-��)���"��uun�A���B�3���v�߆8F �����m�r���W��E&R���kGd�Wķ�'������b��d���,��,X�~��o[��bl���k�֜ҵհ^*����֔u8_�L��]���D7 7��V�FРNj�7K�0��K�"��x�T����؅�P��6cс^�i8�|�_Ф<�� l�-L0��l�?�[�"�)���|�]��e˥�������\:ֹ˴�N�8B��ʢW��i<�DחLq�v���� �#y��,�I��5%K�"A���ڻ��e�&�H9�=�=Yze�~����X݄v���:���OP�9���7�I�L��~61��5-ΡU��<<6�&�(�mF�&r�'g����'�Y ��+�)��s�J�cm2��A�m�m��\M�Aq�~H����v@f�dxna�pY�����࡞ �U�j,�~v9W�ߝîC�G��[�:3�I(d�uq����]��|, EP��������h��u�ڭ}��QD�P�φS�u�.#M�#ZX��(L"�繷���"��TA�\U}̯D�+k��(UUE23��"Ay{SED�_���/0�"��,GN�)\c�FY�)SFY�o�fx�SI���~z0�`���_��}�| tg,�$P���wv���6ޫX���Ջ"���]�����?���vN�hg��]�� �M���:=�+��(�׾gf2��E�t��ɘ�$��+��\�����I�����i@g��4�0+
�io��`������S&����tu�!9�C���&8�w\ҊZ���ȵP9�w���T�#"��&�Vl+ⵙ���R�ǀ;XC�t) ���:��+q�&Ҍ*L�����`ｦZ`��<��jֻ��o�Cq�z/���f�cn���%�\ ��/Ȅ&Q76�m!~~�������[ZCejk��ϣ��w����9RLz�2#HT@n�KĢ�C�<bA`I҄��=�]��n���)��c�.���ͬf'�ɴ��Q����M7Ь=���[�kD����V�`&�����?��Èw��]酘Ԏ�V��K���5Ӗ�{�2J���	�đ ��Ŗ�/M%L���E��n��@M�As�5NɌ�����M���aq@xTPv��pX�<�f��&���C�
��:�.�ٰy���Ko��8O�#�|��qOr�tb` :�CϹqW+t(ù�uD��7R��`��U_=�%��i#�'�BJOD}��p�Z���O��� *�cd�	.W!����3҃��,�48F���-��_�l��H�,��0���?XD�����ccw�[q�J�����a��]ܲ]r�ܼ�(�c�b�C�/0�hQ���T��b#<y��QP���H����Jx<�%Q�bI���P��aڵ'I]9p,���T@��L�΃2����!A^���f�cv@�B�"���^2Z���i��^M48����0V���2�)Qo[��%(a7}��{VLR�/g)���l�rn��6�R"��ƅ4��)�7��
N��Np��(��:{�T~�7M��!�'��ڴ�-�6�%��qy��Sz������4��ѻP@6��-I�ȗ�9��λT�?̛1�A+"�d3�q��gX@/LO��F1$%<
^��*�'�r�^R�eI$w8˻�ʏ%׊�"��JB�8�2X���Q�`lA&�������~��}=��EB'c���a�1�]*��R�^�p�j��`)��H�P�S<;��堬�V��͇Bq�J�z��p���/���H�߮~D�m��	<�LZ�(������nj��>�BuT������a&�M���#��ȝ:.q����b6���e�IM1_�L6Ӵ��[�-EzpaQ�x?ߧ׹%�}��4�!Jj}�ް{�y�y�h[Ct�4C�o��z懭C4=��7�PH�y"�Ӏ��z�*	q_Q�l�(i6?�����j�?���"fC�lg�5(c}<��mSZJ:R|�#<[mAd�K��R�Q�;�68lt�	��G:z!&¢g��s�õ�E�i�.�e,#��Y�)"�`�c���B(;Scwاz��.e���������B�B�Nz����K��ϟ�FqF/l�<������{u���^,�t���v�!���t�r*k`OfM�im�>6�Ţ=ws,r>���J�(�A��IrZB,i��f��4EЫ��[Prb�s�$H�ү�`���_�i��Q�U�(
�y4j����,�F}<���+�ԃ�����'��u��ظ�-�NxȥDF�ޯ]y1���Blk��B��^j��L$n³ �����kR�>�N�븃�ß��K��G&�ߟ��Xx��Z���+h���SbHE8�H���c��m����}��u�#'J��:����j�9a���ɟ�s����.�'M�KHp)��C�z��3��3����}���t`��������yS�3���K@�П6��1�,���\�H"��։͟���l���p\�-��t'&��br��&/�(۸|*E�xX��4��a�B�>��3:*��:���������O�(�3c�F#�������� ��|)-޳�>�(|'~�@�(`�Yv�n�i�;��9B��+�ĝ���q�;?C8� 3  4G�Z�������;{��8�{�ܶ���|$�w�K��R�׿�����	����։���G��:=kԁ�![����`�!T ����[���L���"��=?�xC�h&����e�=6[�$����׃�sOw
H��Vl���LzN��;2T���6L��/�R�1׼��Z�L�g��F�4��%�<��{���XK�kwf�ޜ�73��0�%��n�vf�X�u�xn	��j��`��2)�N� A/D���w�J
95%K$�syWbbz��O�˽�c�@�R�r����Q���M޾���n�ݔ�s�	�'a�V:kϿ�]nT�� �L�c�E�|������D�(Q�}tD���gB1b�����<��X��kK�%�Z&������kJA�w��Y��H���6��X�H�ٺH���N��oĘ�ԃ8�e�ȣ�3����j�	�����<�|����p3��O��o��P����<�#rm�[�K���.���<�A��Έs��DR����b��d�w0-�%.�{H'��x�ϡp�a�d�$�/?��X���6�A<ش�h�p#���Ʊ����v�P�Uɽ�*/p��#��8��w�`)`;̣ҹ�;
�pgmg�[?M �����k�`^=�� �i�� /4��=��X�yN�#�S�̎c
:����f"F�M'��'|����U;�T������ĥ"��QQQ���/H��yWe��i����Y0x�L F�'a�)���C��P'�(�7�AGNSv���:(��x۸Nx4՞fz��on�S�n��~a*W�߻�7����k��{2k����W����T�49(S��z1����Ⱖ6���?{�l>�F�vr���9�*�Z���� +E�h������F̰�w@�l]N`���&YH��q�M�e69,?̈�X�7FJi�?i�
>�)y�����*��U����!�d��z�.�Y�f4��:��
r�}����Z�Đ�M�.�㢽�Z}�%ρV*~ �qW�2�\x�@sdtdQ~�_w�A��hX�I�Wn2��ی�
�ȅ�O��UVei���g�⠊ ���������璵Ԣv�Gc|6鞵Y�l�#
B�k8FC��0����ܾq]9K���I +����$��`�٧�>��J[�l @�Y�v���	k\,$_:�}��5�=>�wz���,n[�$�|ʴΞ���ec?7�B�g�*WN�W�􉆈�[c9����g�&&�mw=H|���M�(@���O�C\uBУR�Y����[�O�UǸ4��Q�I�e��M��#���O����55!e'�aʫ�p�ӁUZ�B�yH��g)+�̍f�[�'r,Nχ{��j�e:�33=~�x X�۽xMt�Z�j�ǘ�q��v��<U3�HˈYlǫ�x
�U�W��Ҟ��W��5� FI <���!�
�|�6���}-@���(��U�w�;uVD�LL{�Ra�~2�NdBa���P�b�b�ݟ)g��%?���=\�f��ˌ��AP�D*j�ߎKPz��AZ�>�Aiʼ�|�e�ʴ��eg���a1;�%V�a��=��4Ѥ�W��;��$�h�T��6T�C��+�3���̢��Q��`������'S O���5���Q�  �ZQ�p�8tT��.�������p.�y�����ҵ� �8�?^I������KX�<K}L�J���|3���F�+�(��ϝ�]��w�6s�J���U���n�(�v�� OD�m�/�I*أΰ$b�dM� ƣi�10"���jT�;��V%�n��o߽IhQP9��𭏐.��礌Hu iw�
$,1��~�G()���F�Jྊs�W�կ� � �Mn^տ$���}��/�WjE[u�����z$����a�T��33�I�F���k�`�PVF��m�,S�L��s7���brU�.�R���a���@d?��2<W��(�/�茇��EG	�OR����9�`1������q�'��p�[|��/���U���:�W�ٷ`�v�:Ne?��I������;::Y�b"\�s�I���A��
��]����C��C)$H���]�ږ�q��ل����3�	�}��E1�Q�b�r�w� txҦ!G�G~���(�MD�,�ܧ;aMBZ=��q�5;�I�h��̀o�_�����ڹH�v�h#���� މ���6"�VJJ ��E�%���s1?R;o����%Ӟqk�ҵ��/�
4R*�����-H�2��<�N�H��N6I<c����֐>]aDk���@U�b�_Zc=ŵ����Ս�{��E��P�:He@��\���>U���`���3�򺣋��8�l�F �׮�[Ϯ���t���D9W&h=��1�H�[�b���	R���!Q�;m�����^�پ�'�u:l�Z�:Äm~&Z��@��;��<N���Q�Y%@M�s%����g�r�QC �I[�Y�����>�� �j��;s�Ή���58m�&a&�"E�&.R,�aE��V�Z-���Ì�t3�������oOܨɊN�}�#��3�������@��j�+W���[�����<��v����L����ߡa��0n!��җ������$��Y�F�o��<*AGhFW��`�>���B�V_%�M�9Gq��$&��AX:��m:�����k��C0H�i��<1P�q�4Q�kR��Q��EP,�V����	cc��c����oi���~�S��&AJ�������	���}vt�%r^%:���g:�`^�3���J��GaѲ�`A�> #-�Ab}��d�/���_8WA6!�HǷ9ׅ��
R�!1�\k��^H�6�R݄�!lL\�i�b(�1\��^˾5��q3o?]�`��ɪ��W�n���8�ROo��/��/��6��`"�g</̽ES<b[J���v^��ٙ"���,����:��ۖ�A�K.lO�Q(�-�x������o��ݬ]̡e�P�\�j7�aP9}�,@D��d@_���p�P�9ʓj�7�]��Q�K�z�+d�o��ռ�Z�Pn��O�e��&��,�r�_�d�d?E��B���ll*p��mQfϸd���Q�2�5r[�I�iZ�W�H�V7���É�쁯�Y�#*!�+ǥA�_�I�]��c��L�} b�I��;D)YI�T<��oh�W�b�ơ�G�L��yJ������_t� ���9��{-L%T3s�%��7���3�����|����(��m���#B�݇�+����SаKi�q��T!ۋ��_,�D�{y�f
����q9sAm�K�P<��٪'��Rv�KUm�T��bTxX��UvuŽ�J/�r��翅���]���+�h�e�g+��h�z����b�պ��$�F-i���k9#(Z�Elf��|§���yMU8B�e��! *��\�����t#��Eu�bĝ��M�/�[
�Dɕ+�1�W�e_E)9Q5���7+�kW�S�M_��U���(b�[�@`o~�/k��3�ٰW��*D���.ys`�TQҫh�Lfh ��y��X��/~�v?9_����>����i<����j0[�;%|h٫d`v����,�q�2;�zf�qq�<|΁��"�lw9��*2d�Uo�P#M�Σ=�F�^���F�+����.�O:v�6���Ȗyd�	\q�+]!O� D�8_����Gu����[�_#_ÕmبW{�)�bc[\ ����'?k�B�t�¾���1�Q����{���[F�+���L�!vH$�0Īv`l~��\e�7��~Ɉ���'�#��>�CX���D�u�
n���^9�lnL�o�c���6��CU�Q�Y���I6�X�/����S/�U���x�`���� �Μ�0Z5}�cx�L�������_�]� �T�ۧ �	���*��3�p�%L�%���-ᛚ��Z�ma��|c���]ؿ`�櫦^�-7���,��@vox�u�^�n�p�Og*#����B$-BY&s7W.��)p�|�?��1��H 	���_8+cA�z��v�`]nw�lB|���VKQ��<)�|OAx��H׀�E���K��w��c���w)�3��	�����8I������_��'��=èw��B��S
-���^_�_7�R�^�I��F�;�ĝW=��c	�ޘ�+a��^)�G�ֆ��y�`ڿ�5��u��c�M�=���lpo�>A%N��+1�w�P4wViqb��SFCЊv�դh�y����G��h-�������u�48��#��9�`f�������b_�#G��LT���04!�55(�#=�)�p�����z�P���5!;�k�91��O:�r�A][W���t4Owp����֘E����͈�-������Z^���������@N���a�9��8w�0^@~�����=�u��j��tĹS�pz�k�{�J��]�볢�+�;@P�|�._k��A�]	-n �d�1�d��q���/D�[f.�@��w͢m��A�(�Zİޤ�BX����;��W���/BpfsS���6D��n�ð�l7�z��(�UR��<������?�*u�����+z� �~(���;����^�Ne@�%���p����R_٤�R�Q�w4�a@�IA=We��E�-kt������9N4�Bs��b3�"�0����p-kA�sl�a,_g/2N˛���U�:/^y��eW�5�
83�Z�lr�|�B�iv��Ut9�pP8�;!yX�ݞ�D2T�CU&�%>�1�����27Hi	abͻ�b�83������b��q3� �2�w���r�}�t�LZ1�i}���m��Nât�wp���o a/ڰ�qrs��W`��&�ޮ׶���ғ/Nq%�?��.��j��Ena�a|������v����	��ˌ
2^�]ǐ�e1H��3t�"�Dj!�JxR^Y�4@��air��a��5�B�B�lm�̟��N���,�f�(Nl�;�sQ���6X\'̯�`O�xW�N!���}�Ꟗ��V����_	#3�*!�J�A���a^�����HF����{���P�oh�kuf�*ʹ�=8�9�*�,��3�48��#稈��/�..�9���5��?
�����wok!O���Q�i�E�G��|eK���U�R4��Z���"��;���_��|��@�b^y���t�`�%�D쓖zdi�+�YeS/�CL�s�n��j	!jd�����?���m>���Ćީ'	�nˊ�g�-xf��W��&]�q�3u�'[�����E��whm@&*+��<ƒW>;�M������t7�أU�sk��,�g��b�($I>��C��AC�vm#1���T�,�>�y�A�)�u�B�cL�|�~�bd{�g��=R+<����c�fbX�%Y�I4�γɒ�����o���ݜ��vHI�o��-��{�`��g*]�IA�^��P�~�]�!W�[����k�ޠa�Y 9ZF�`<�w�c��u�w��\@T��h&��w�"[)�����-�l ��d�k�|��E����٫�et��I�gxH1����|F[��$��r�7�
��"l���H�	7%�gg�'z�9XcJ�ǎa��/ m�k�7e��N4���/��+�U���>�P��k31^���� �!��1����V�EH�Jn�Bqx��Gw��
��V!`9 ��t..�+>��������H�~*4�1i�-�&�w��Ha� ��m�il�g��)�u)�
��� $%�{C�u�]�CWL�PC�����ǔ�i�;�5#��� ��͇�2��[��C#@�ٚd�ЄX��&;�6+K/�O8m���YzF�!ia��IJ��]��qKWX�s�%�%���%r�cB���e���/v�cC�ps?�7�Ȕ��@ ��~��9���Qfwe���^��:�՛z|�?ˌ��G�$Ky�\�b��r��*����hTN��?]*��42��7��r؍;�Ћ���7���� Hs�"FQ֗v�7�	�F�KGI�S[�𱆿q�v�u�ty���Iv�/
��� L�[��c.�zkQ�A'��?�Χ��~K9�i>�^�h�S��`�DyI�O�pU3�3���3�B��0��ړ��}׊\E����h8�߀?��}�/���DB��"��k	����}|B�l�T.!o� *0𾋅[�£�WS�3@�rKm��	)��}�祩-x>[ݿ@A��pEw1>��`����w����좾e��
\�e&��?��ވ�}�2@�'���dHd�5��H|�A�haz���Jʾ�Q}{�#�qV�c �ڞ�'��f��;�bT��M�ApC��Џ�
MBZ������y�,�+����Jy����]J��b7���������U�d��֓X��k����bq����h�+��,N����o���͍�k����N���ڇ��k|G[x�|�jt1�v\�Aͦ��&XP)3S�x!��`	�F�V3��ŏ\a���;�˿w޼b���I��)��XI�jmv��h�F�%�.�R�i�S����q���:P�ܥ�"�� ��$�|��%w��|�L �����ɟ�^�ۈ�����8������24�]
ř� ���h�^����7�r�?Rn.�'+޺;n��d=9%f����Zʂ�I}��YE�MY0�i���{(R@�d
0du+����Ӳ��1c�R�X�Ɋ�VAd��
��n��c��ꗣ	̈���F�o�6w�.�������
l`�����Z� c�|o�M6A+��^U)Nቆ��P=Q0���@��gf�A���"��1��ѭ���Oz��y�`��6t��<_�i���aZ���������%��|�m9��sD��3��}p�Ґ�@eC�� S +��ѧ�	fô�������g`L���E,�|sʀ��h����nݖǑ�Y�k�:�>�v��7Y7�$��
j4˕*�(�dl�2$����%,p�#	/:-BB���tr����GL
�(�)x}뜞����<v�K��D���w�hg�0�E$�Iᔦ�o�M����P5P"?;�r��F���5/)tX�`��M֖#/�YOk8+1 ��v�E3��3�4�O���k^��(?�B{�K�n�Y�L���}��YɻHO��/]�Z�z�=�<0���K!H�Z4�L��t��qb�/�:>D2��*���_1YG��}�z��~b^[GdX9�� h�ߓ�)�r+<	�����!���*�J�N��<p-����I���9I�]�]�1�ɏ�*L�����mO��*D�A�fPSH�WP!rgɝ����]/�H��?|�=�"��l�"���fZ-�"d�D{�>Ur_�,�b����gl)�/Q�v��<+b��]��B�L�"��ɮ?�����A@��~u�螐눉��&Ni#�� ��B� �h��O9V����Q��>l�;s�x��$�� zf�EH�l!�n�Gb6�-�J��`1��S�vz�(SO������K;xDp�M�G���gi�&��jۢa|긪�C�͠F�t<b�:��s��٧��<Gi����c�*�4d�Q�=e�3�~BbiN��#���.���E�'��Z;;[3�$�V�Ͷ.x�d��W���X��X�������y�A�"�F�N» ��:C~Ceo�`��~f��kz�Nz�w�K�����)Z\ճL��z��<}����1�l���P��yۧU���ɖ�&J�}{#7�Ja�V��N[^qݮ�l�ߪ��aȃ���&"���!���FI~����W)��я\�5{�T�+�N`jh!��[��&�J�e.����g.���hV/�أ6�� �Kry�y�`x�=�����Ÿ]b!i�TA4��m�H��H;�;�1�?�޿/o�{Z-S���}�l�t�w���2c"����S2��}��~w�*��W�S�ޓ�hg-6�0e�]����GH�ѲF��T3V<l
��a�}��f?��f�:��塭JD=�����"�4F�@�'��2OS���V�s�tqQ׃��.*_G�\����!���cİ�i��
F���V�x�qT,8iF�v.��)���� =��`UR��?�G�H�M��DϮX~Q��ֱe��kjc��~��E:���w7W�G�R<�p��m���s42�@�4V @;���������)�0z̜���S�$ȋ|��[ �4�m�(��k��/��c릥,��U0s���A���ۆ3v�ˌ�nm�����>ງ3R\�c�2&O�_�������|���d|թr5=t�Q���}�5�-�;���b�3��̓3)�������	\~@���e�s�xA0����@�� ..4T��1rt+��ɕ���I�8PE-чi�ݘ�4�-Ƈ�֋F��������ſ�N�x�?I��1���q���5%9b7��ZO?�d��:&п�0.�ӛ"���C�۞�{�]�P�+�.���Lo�uQASO�몟0���X/�cΆ�C����若v��{AV��RY�C''�==;u���>����%�0�X�E����h���mX�e]��B�)NM~����mD�#�L�G��"�T0�W,��'�'Pxw99�α��BcŇ��B�E�)H�?��+�-�6�)��q��P�r{�p���ǄV��lP���5���ܼ�W��o!_���ޒ�lm-���о,9�؏�w��Ǥ���\d�J�� _�i�aG78|���j7��SL��)Sw@ ��&�5����t���
���<�e�aފ��u�cn�28Y���2����tu0���b�!I�b̦[W4�H����@d�P��\9�e>թ�%��=�pp�r9����6�|_^�V�f�,F�vL1���,�"���Dy7G��m{�ϯ��S��z~�ߥ��ɤ�g��~�>6�2����>���O�-��<�K_�0+5�V��v����ت�]5�m܈�F����#W߸N���֣�-ze�l"Ɇ^��}7b*���GK����L�[e�R���.�̸-�aW@�Dd߸�x��]M�6���j����c2y"���8�W�����;�c���.���e�Ś�_��Jҷ^�.���`���G����8_3�s��N����$*w)�0V���0�O#�=>�c�<�ټ�)��z����Ůվed��ꨐ�
�LM�!�����0�EՑ��%��U��RB��%Գ�,������~��!uc��9h��1�nF@P�v@t�ѩ�^h��d���,%��k<i�w�u����fw]tU�$�"c�ϭ�f>����%�ih~Q�E
m>����ʤA�+k�bՠ5���̀�YY=��lw���1��PGF�A;PH�-U ����	nH�S���={���D&k(mG�,��8B��+H�=VV�&gfs�7��<<�lO�_Kc�G_y ���&��UEw�fK����E�HS�
���Wv\e��G��o=�hj��C�S�V��Qw,���� �S��a�6��A(�0�l��Xs�0Lh$]`Ν���������T�����j`�x�=;/]���RW�� �����{aA�j`w��;U�_��֭\��m"]��n��fy�P_O ƕ�N���d�ɹ1
&��ɗɟ�?����\/p�%ӦHY�n�ā��b����a- |���)���ѫ��F\�I],�h�Lr+����1�8�aLB%輂r.]倞JE$�C`�ܾ^��I$�$�q�-�h��4c��V��l�sJ�}dA ����JM�$�8�����%�U.����%∁s鉀�v��S�vi��3�@m2~[z�a����E<��ǦWq�M���7�`��T�8��;��ai����|�KLq��GN��6Lr5z�8}�� DA����aO"ĵ!!�g9�-�a����UTʁkx\���>�Dd�Ю�L�}n,�r�hʦ,�X'#�O�T,�Y��E�_��r�rOM?h%@ֲ�)��c('��7�N])�@02��N�f��w[S(�gF���׾l���!?*8 �Q�H��k���e�%�`�&�DӚ�\A���M�� �R��/#3#�����:P�&�_���>��7/R:�ev��� ,�8\�t���1WK��(}8�T��KQKcuG~�8������h���FI^R���K�җ�E�Z~��,+/���C;��Xz�֔:��
�$8��&���2A&K��f;�S
��u��=8�Zy�#]���*o}p�P~9EK�@1�v��P���El�?F���^�e���\��*N��ƫ.�t.y�XS�Z�Ɠ#��t��!nQ�_�-��c)���9A�!����[����{����D]��'�{K0n�-���~�!��\0��D�IZ��J��"�YSD�V�����Ob�#�QA0،�l�R�#y$�@9!n���`����o!&���7nt�^SˆQ��	�ΗM!���>��O�_]�I��^m��j� F�N���>1v���<���\����t|1��m�F��qo�|�n:W���w|6�z�c���?1��H��N�������,H�o�U{�B��8�����,�̦���`�8)N�]r��q��A��I��o�A��!{cD�4 ����������	���퉐G0Y|�ƞ�����%�!6�*����\������q�N�@�ڍ��h㖟�!�����3
*�����k&*����"�5axJAр.�^�<���ר�-�,��A1R�]Q�Z�o��10�����#Wrj����^��T��|����?%f���o�	�n�|X�H{�Qm�����)��oe�(� (��A�we��֗|�E�^ʉ�^V@���
�(V��1]�
�DŸ)�͗V��+"��U���i�%$4�)�
�ɮ}�^`�l��h�	�o���Q&�w��Z�i�V���b�B�Dd"%5r��v��ħ�E�3P���k��T��z�l1E�_;ɿA��#�r�& �$��e�C��i6@���ڻN&��� ��;�nɢ@1S��I|M:�çNa��fƫ���rfX2�<�m�j�UJ�j#�cZ"רg����~�$�r�k�\���O� ��ef����`�}4ݴI�r�%�p���$����aۧ"E���J���-_cY��J��a3�C]�2�"�8/��S�k��z3M�h�bT�IDx	����f��k��[�����<և�q(n�\S9N��Y�Κ�F8ٺ/���������T���2k�L�ݡ�OWe��:�œ����s������U� ��d`���B}��ŷ��1���-j(pAd�+���k�6L^��#�ԭ=d�3����B��0��7��^~�x��0o�hGDƍM�����_�2�w�����`���<���R���3�G�ݱ�0��Lm+�2<�
�*���Tx�I���P��p��Eª��r�9���<C%�R�2����ŋ�r��a�'7�)��{��;zQ=irR�m�ids�P.�H1"�W��V��Hr��Ȉ���!�PD�����7�]� 8���&��7���\��2<ؖ���������7Au:�xi�᪋��k
�yX}����,�Ӻ���L�V���=��_��wl�ׄ��@��[�G�'r(�E��aݍC��h"ZG/n!і����(Ԭ��~WzV�����e��%��UM��MT��ć�P�>�r�7��-lQs�//e÷v�SA�ER��s`�)����Ù���._�R�L97Ěi^�-Wdh�T (Y'�����,t���ƥ��lm�0ux~�<�T�⭸*, ����FcmY��M��T��g��t;K'fk]A��d����)6)=��`OH�7��yh��v�����3���/�|���*�W�L�q��w�� pRA���c&��A�Yj�ZNq\%;Q�^����'���+��������|wjjb��	�b�OJ��wW���:��PA�3������AJ�@<��+�R;5w<��5�|�
�I^h'��p�2y�K�G���]�mZ;�3sR|�T>:a�_�����-z��c=ZT��joT��'ލ�ZFn�ͣ;� �&=�m����*a��?��nBؠ�4�}��@����
�qi>D6!�V�;U��Iol��{�/�Hﭗ:m#fB��������2>�;Al��������[-�%:�SJojimpNZ]��QvbT:��mX��z]Ο��H['4�+G�C3c�pb�6���w�%�\�L���~݊$B~���+G��9�y�}�l��MઔCZ�f-5s0�͹R8�
�3B�qv�V��2I�K�W��
h@��-P�� sq0��6{GT췬G�3�%�2f7�)G�ԙ�&��,m�-X�u�	%�<6@f̐�X_P��5Y6;�ťy�rQ�����y���?#�7��	Ɨ�c���,�����+Wi$�U�Ƅ�Ye�ʅ:�I�s��I�D�t�p��5ꧢ*:
�>48�|s��֨��~���D�G�_�6Vv�I���!E�,��M��L<��2�=��G�����bM5z�q� g�ґ?M��K�ɦ��N�Ƽ8�`#���.�|q����X�S�]_!�/�?E�RG�4ߝ.�ϬK_h5��@�J	��ưG*��4��$�� �M^��/�Y���Ԣ:fD��y�|mE/P±j/$"C$�B�:�	�> �p!�p�T5I���^U��,������!�_Ȇ\<��7�Q��d
rD|���(�ۯ��w=˷��y�I��d��x8$��-��ͭM���#Q���6������9��ыc���f�^�?T�z���|�:�s�6�<5g��h�\䶦NnS�V��(�Wx]�0C�|����lb�s�xS�f� ����ZL�Qk)��)���Y!���1e��@9��.H������ �, D��U��I<� ��Fv���_��|�+@5����x��,�ü�j,n��}��ȱ8z4IHR����AyC��s�@�G�v�Ҁk�NV�kI�갭w�p�|��e�;}I�S�<�F���Z��Q�*���NDEo�h��10���E�n��'���!����#� �%�L�$p[Hj�5��C^ .��	f�+_�(wO�}�n�b�v�>�*��o���p�]����F,n�w���n{����PwQ�-�O�e3e�gH�դ,¦i�)	�<��*�yP���I>���Ꞹ �[�����%�?����<޶��BP��Uo����O/�փ��jM}5-Wl�k��D����*�8w%�����m��;��Ȱn��Q�W�8�T2}!pY뮡�DE]}��:՝Φ�`�I��:��zM햡>�w�/I�go�I��r<�4�Q�Y �x8��/�����Ł���p	�cB/6�+�
?M�E&��sY$e���ڤ����!y��#(a��bw������j�)g�ƺ��Jv:(��[^^�mƙ��yr��Bx�K@�.O�+���%OzؼDQ������f��u����W<��ҕ\�����tz�b��u���F��o��M�_ev�hp��9K��_x�6j���l�8�q�"˶{�:���n��� ?�iU��߾���+Sq�����!��tQD��c6ܛ���8��Hn���*���7Y�R\M#i+�I�C�M��p9���{n=\&�����'5�A��h�&
�W\����3�{�)D�J�|_��t;9�1,6��#W ��� Y/�~�ԫ���	'�S�%m9n���6��# ��׍I(��VOZQ�_�����Y�+8ķ����vy��M�V?��Lm�&k =n�[���:�u�Dv4�Bo�[��� w�i�Q-�e��͌a[�+�j�H����\,�%3�e��i]H9}o]�N�my���V��X�&����Z�9��@�SI:#+U%��7������#|Yf8���0p�o �m��yW�S�e���'sw�<]���[h}7�b偧��z�<V�(�)R�aXs�y� Ioښq�F��Nm�wÃ�_W,����V`�rn��
��f�����C�������;� �%���u�,���+���84f������T@`o��R���>\�f�8O	�i������Sp��E5|e���v���_{$��Q������&:��ٶ�ߺ'H���r���H�2�]s���f5%�.>_W5���5,+&#�ʋ�����S���(9�$�$�Q%zt~x��Z!b �KE?8����U,,��Ty��cV$3-���[��i�?;l&�{��s
�^�#�o�B���bE�|+���Ϩ"U:�D�'kW>�;�Kqܲ�/���o�r��Ș�]�S%Rv`@�)OP��=�z����C7U���b���T.IP�	q	�ט�o,i�/S��N����U��B~S�/�.�F��$�a�����e��L����G*�ǭĿ`�e�P��O;�w�AB�Ԅ��A����3A��\W�G�q��X+駺3�Żh�Yu�����<0�]gg{��e�S��!9!C�6F�f�����,QR7�A��ꢑMܡ�a�mE�J �"0��As�4�ǌ�Zؗ����r��Bt��>�z��ߥ׶ �`#�'L�2I.P
�۽�#q ���#&W�Tǿ��5^��_K�g�}�e�� M�9abʊ4�4�ݭ��1�������xD[!̦y�������@�F�?��rx0_ު�lg&lt�y�v1E`}ҙ�VJ��,q��[��'��c}ܮr�̼s�*�\L�+��ڙ!���O1���'�G{��9k7�V��;8��QƮ��XM��)"m����\dd(:�+[)@Z7)[ෆ Ϡ�|�n[��:�H��x#v)��e�+��z���H�U�I獕'�	�䎐S����Վ 2����9*m�]a���W�]�d->x [�2#L����[X��h�?���;mS�O\Ѻ��Ӂ��bn"�W�I)~��s(*A�~y�}���ϖ�c�L��D���;�������h<h
;�ܣ�+Q�>��$���A9a�!���L�����!��o-q{0�as�C������D�����f>���s�!�uc䇀Q=��"�X-�Q�gOқO�ѽO2qC�V�U=��?ȃ�_�ڗ�+�ϼr�_@%Pه̓�(��1�G���\����PD��mڀN�<���P��t�#�d�ԗ������K] P�[�I�2':[D���*#�eR��N�)
���)!�J4�L ���jh�mlR���T�A�)
ɀ>^|#ﾡqÏ�\�$c������rm�^b%S�ЅL��rV`9��F#+9q2��/�L��n�ROs6��a��>��L[�5{��q,�No�B$:'[��a���M���bEwb�͏]��6B�c�Rnm��T΀�A��x��j�2Z͝�t��u����)$��=K3��e�B�vr�C�H����xxA���a����p��w<2���~�<���r�����U��,�1论��a`������a[�n��,hyH8�	�ܧ�]���3�c�
 m���݇�	g�I%�Y�s���U��MC�Uz�oQx���6�<{)�BEX��~ &�����R/𭛬�-�~X�C��x�0U����i�0��UO����.�� �f���@Y��\1�����!�_q�0�Y���� �F�bh��'%G��c+ީ���D�mɃ�=���Q�]�.�%�2o�?oB��2�i���T�Ǆw9���Q�$#��u�i��U��1 �[���ǣ�g���аP���֧��ӗԞ�J�����C���NY���S�G�4l*�	��I�T��L��jѸ�V^vz1R�]G^K9��n�d˩j$�r��xYw���\��|���O�h?�Z��E�����O+�5��.:�o��w{wP����'MW��K��o�*����d�R�$��,�k3Ε�`!j��r��7�r������W"��ނ��_�/a�lH.�aæ��h�˔��?ם}"��<�?�@��O[5� �Zuod�}+��Qĥ���$�Ts�v��b��sU}�3��l�4	��j���A�7��ۯ�
1��2���
���݈�$�!'����q����ȭ
��E�0�ޘ��k:��V���k�{�6z��?�C�v6�Y������kϲ;VѴ�.��7��v�jItL4cK��s	0c��#�>?t�������mD����Y%RalhL�<q�P_O�/|x�`"����V����ű|`����_v�MC>i��C��)�`�=,ġ��<r� O5'�7�y��*���-nߟ� �>5�¹��k2Vψ�ZET*2�$z묒�Q&N݈C�杩̗��?�j���K$z��2�1��"�^�_O@��gᄌ��}T%��^���}	��pbr ���KN��Ә�A���v)E3E��>���m�bM�Y�'V���K
h�&+�r��V.�[��A�Y��C<I^�MfṿK㈷��%�G�[ʄm��ns*B0>FW'�V���F�4���=�B����e����T����tL��%��u��;�u��ͩ|�5�ݩ��:H����-
����]��>K7WD[>hR�T<��4O~��q���-j���Ƀ�\���GO{�W�M�oҴT|�[�<5�P4�i�cr�H��1)p�$b�Ƈ�ވ��k��¿�5管�^KW/��lu=[D���CZ������)F��?�v%�<�͆���A��4m�x�Xl�_�t�@�Zޞ|@�ݬ�<4�D��d���v�`4P��:i�6�]U�݆a'DlVq��U�84V���8���[ҖrI�n��X�� �'U�D�EO�\?ÎD�Ǜ2�;�W��Ќ�y k�R�#��҅lH�%_�؏`�����1��1���{�q[pj�	sx�4Z���!�ul6ۀ.,K �[��n������nn�>�6*X)�`L(����MZ���֡I���%6i��?�x�W^[���"�U�V�-=�zK��%����v�we�=[E�O-�MF̫�X���ҹ��RZ'�̋S5���o���nG����R��}���}̻�2�J�J�.0ߚ>���'�8@nQU?0'/��:��`���M�.O�Wi���ت!DAl�D"���l��7͏���y��\s�?U/��r*;�\ ���^��o� !�����E�Æ���%��K�Ǜ�ޤZ��EZ�0Q������H��V�:�RO��a�/L���Us��7(���?	�nL]���M�P�\�R���oF]@�L���%��OWܵ�;k/���Jy<��� Dy�G���ǟ��_.�0\�۫��,໊�*e�nj�)K!�]��.�f���(K%/l
(�SX1���,M(OԽ�L͢�y�W��9_Tʾ��Y�t�_�I� -uD�.b��^ޘC�i�W�-�k��H�.xM|m@�R�f��	�� �Ve��Iղ�Ȍ8|��A��K�v�FD=Os%��Ԟ������y���[�ZU���3��)�f����d�k�}鸴�ϴ����q��ƽ�A�YdP��ʜ�^
o���dL��^e23	r�[�_?�y�>���Ɲ���f:���*s.p=W�Mk�g'����o�U���*�}XLo�93��u,B��� ���4<���n�7�Kb0���h���v�+2)\�B��JLF6WE������A��_;,��
}~r�z������r�FӭQ{��v��wC����T(�w���9!n0$ٵ��.���Nmci�HF�����W�ψc�#��l�G�š��}$��-�uo�����>�Q¨�*=�������-`��sh�K2^\�ٺc ��.���:�&���?�{����t-��ϳ_��������ļa�N�3��wU}+��~�ռX� ��?�b�^<\q��%f��$E�Պ'2v�7f�[����C�saNe��5���~f����K���@���?���ä��T�@�Ac��&�ʮ�n�r8erf���j'YR{�Eٌ�?:³y�Y�H/iV7��'~x���0W�����&������UE��^lg��G���.භ�0e� �T,R����E'R�vI���5G���y�����!b3��=�aH��V�W���Qn�]<^�IƇ?J�u4��QZ]1X
� o��bME�_T>�����Y�����E��k����n2zŮOչ���	��@�1e�����!3o.��]���^�v�3�e�Y!q{y�>�>��O
{��E�x߯/�y�Ŝe�]��|O�a����h��A8^6�\0Ks/�����n�t��+�$�;p/(+Uc}� [瀗W3.�_�7��l�6����K���?�&�^�e��4Jڷ5�e�����E'CޭWim���44�gs�屡&Tm�HV�/H'���vy{钍t�K�$�������"fZ\��ߨv��GBrN:'-^(h̩�&[��>��E�>�����X�8�p2i�ӝ�|��(Iɍ��V���89�mD�y��9f��­9��}�Ư�Zl�4�R�~��H{�]wX�Xe'Is���*5�V_;Gq� ؅�\bR��]u�h��=XW���/�?�O���=���D�y��2n���"�]/���Si�r���̰�R�b|�����)��C��� ���U���)��T�(���*ezu�-��0o��~c�QB�3t�a���ۯٻ�񔖋��U�����,@'��J�}:���!�"�'����J�����33�Xm�~�){Ds� �ݺ�+LU�g��߹�/�#��b�UW��~�w�!5���Un�t-&i��wO��X!��#ȷ�;��p�c
�`e�x.͡�57�h(9CB0�]�-.�E��n.R j������Z�+��_?��6 MH�^��
s��G�s�poCM�!������N\Z(��.�#k G��z:�Ҵ�+�c���?K��0nV���5N��:+?�t(
7I+n�4@�?�iGǿ��`��>��tWx@#Ms��D��`aX�}V�&
�Ȱ���H|f�9��;�)F�W�xQv�����"��tt�+	���&����D؟+ɝ�ٹ��c���9�U���N��H���c���a���^�uY��6� ���S�����kl/.�ۭ����l�:�l��m����].��t-�ļ��yJ����=����Ӝ�D}�U6�P_p����4Kѣz����0�cN_���	�L�2ǅ��_�J����E����5��_;�<����5��mJx�e�G�򙶱���؎I�N�ȼ1��Gd�5���|��b�/���%�D}/hnZL��8L���(��u3�.f7y��ӣ�`���D��mN�IU�����ő�ԙӑ�V�P;\���X�D+����e���~��1G}e��+}0��c��ҢJ\�7�  �gS��>���q4��^�����Ahh����[p�.O�h���<:����Zf?���8%��eá�T^�`b{�.)�p�����I� ���w���Ցߪ/!z}ZA�z���B�1��vo�&hNN���l��ly�£C����n�b�"9�]BxVQ�����\PC��EB�VQA�qx�!]�6j����5��_r(n}}Q�_��Ԟ.�>��k��wO:����(?}��P<�iXxg�Q�6'DVfl!lh�QͱdE�h=I�?ڧa�[ٸ���4�E�E���Y�;�fF�p�"�QGͺZ-��o�h���p�yԟ[�Ɋ�����>��I���P'U�u�ځ%�o�Ŗ��8Y�y����F� V7s�Fy�]����҈�TI�9��3��G��|����[������-�a"2|���=_�<cY��T�!�&��s֋i�`����cj���΁�b�nxՖW�v���^�w-pqJ����8;�*���I⤒�5��gl�=-��^����5�J��D���yu!�l�UA݈��p�X1#��ҫ7����9�%�`�Գju�Ixh@���=1Ν�ۉ���f����a�@fɄ�H�v\�[�8�gdo� lͲ�;GK7:���ζ���P^�1Ӿ�j�,&ޚ�B��Z�<5��!����ʤ�/q��ۢ1�YCZ��}r�U����8t�R��@�(�"2J��Zt��spy�D���S�\��xdƟ_�u1@�����Ty����d�ws��Q�R�<�bJ���dH"��GU�hP-�"��W.��$ӭ�|2�-�U�9W)_�??��k�y��Ү�G�����
K��.����}�e�������,�e������52���6F�	�KU��'�~j�{��4DҝL����^�l_A�/=.�U�Q[�玹a�f�h�=��������y�\��~���?�ڝ�>(�ҍ*�����q��p"�`nΊ�M��e��a�<��A�b��sV�'3�� +?��=� ��!�`��Ʋ�3��gt�L���`K�0,�t���c�IJ��D�\z�1�tq?tlUI��.�@�=�~,t��@R����<P�n�"��i]�H�t�>��C'o���$��ۥ�z>[RK�R�̾����o�aA��Dz���rS��n���H7����zT#0yI�����Δ�,}�[��䔑�޴�}]kYZ����Ϧ5u�
It45fk"ů\uF���m�|cN����FO̀��fH�A��
�E
І�%bR $�ǰ�AA

�#�fw�hާ��vU�N�#.\�,�.�l~���B�,���s¢|�J�8s��؅#��zi� D'Zo?ok�w&?p������W���?�s�G�^�T�30 R� C"�wB�����^~����+�I���Ik4��C�qW��h�?~�^g��j��C4����7�}�x�Jo���P�HZQAuw�{O2f�-+z�x���q����ZtI;�=DuV3	�U~]�^.�VNz�
��#yWn���
१������0G�"
�<Z_���uV&����PN<����@'�$��9̣�F�*�P�-�*%3+��X�F�G-����_f����-w�:�H��p��Ig�4٭��N�ϩ}d�]�	�o> jj
�"���ȋ�L_~����Ol�Q ���
_�
��Z��Kf[�%jB���L����O��6���橐��%@�4�WW�I�(�o�<� [N�i�}Πt�\�.�5���Ec��q�O!�S��H�Ĵb�������HP�#\���w�s���`�P��r
�C#�l���}�d�m�fؼ�$�qL����r���S��庼�HM�q1�֣Ԝv�
٨�j���F��?�C�2�<
c��7(�Im��0>{V%��UJU�B>'�Rs�!-u�kc ��4�|�8�\�X��ttR6�6k�#I�"uIi�(E�4��(A�fU@0̸��Zm<k�P~j���N�^�vW�K�A�N���1K�� �9�@��ǻ_��TyͲ�f�p0��i�:��g��	.?N�%�<�?�^	���r\"�>���p���7pP����.$\`��hlb�]'8m�0�Ez���k8�`KZ{�a�&q���I�10WZ�'�z��O�hU�W.�%��d�e��7�hr*O����yin��J��~CH�*n������p!O8%�r�_���Z�c��l]jd6,��-��D��dd�<o����m�e���|�!��JF�q�)��!�XT�\~fl*��"Da�h��r_��A@�1�b��ʝ����,����(S��� �Do��4i��@��/ڼBk�d�Y�ܲY�h+E�M>��S�9V�ԗ�/���9Nʞ�Rd-.#�|����`i������`�p���7�r�#�>{c�xt�'��y�]p|"cj6	R����E1ͥ�O� �:\u%��!�GOĐU[�3R��3X�$����c��|�s�[���Ԅ҄���mA������>z�VfbT��t�mF��@�|�/ڼ�iѕ̙6�C���AH�m�e�9�Jw Y'��Y�ć�^�Z5����T+�4��+Ɩ�ɖ�ӇL��u�wЕ�ZA��S��Zx1�?d�?��T�Wi���}ui�FHR~��r��A��B�*D�;��򏁋���W�g��-U�BG�wv���`��gڂ7���8B3��p������V%/���w�y���q
4?f�Mǜ�=3T�7�O��+lZ9;L��������[��*�����o�^tUt>63����c,@����Y�Z���nv*g��+��p��UE�" ���ߋ"]�p|�\:U��ȴ�I�v]�N�|��,����8�i'�����'�?� ���M\���n��n�����j� ��:��D�M�ݐQ��VX�nM���k��\��oU��$�b�gȤ������������NԱD��mW<�n0���蟔�%o7u�k�c�*��?(��QN��dd��������"s<�خ<«7H<� �_N�4�U�2��M� �O�m�r���X��>�91�W�٣�9��zKG���ZK���t���H0#��ͯ��9�7���j3U�����������͔"k%!���� �et5�,D��9��,��˶K ����Ђt�f��� ��c}�K��q.�I�<�z�����݄�"�=�|�ݾ0�&O��\Ї�9L)'���C'�6п (��Ĕ����3'Upz.2�O��R�#�jwΑni��e�h���<d2���~j��h�8u��Փ��z~)����T�-7�)jrz�#޿����Rve�#�[}���[��R1��݆x�v�~iJO�l��n�վ�#�ϑf��D ��Uh��c;4�����#���Y/��e-�8��9����5�a�`�xKn�mn:MY��\8vM��[5u�,(�J�N�j���%m�'2��a߶�oњ�kic��67-�������rY���/��?��i147��?�/F��i�P�OY��/� ���B�42�d˧Ag�;h-&1��"6/�O�]�l��ɟ_"hh�o�QG�*J���2�(j���X�BR�
7�.��
Yy��XPr��cNA0��
����3��ٳ��%�Yx��\��|��QL\�|p��w"L5�������D�>��>���mL�V�P�M &��Q�E!��|Q�Ha'��~$��B[G�ۍB�q��*����/P�ܿ煫b�m��ӷ,�~�%��P(0/i��Ns�rB���2�<�l��s��d�liN�B�&^@@T�dB*���v��Y��4(���&��u��"�^(�ϣ�;�*�4�y8~�� �=%t\���,���nB���i�n�G����l�f�b����G�}��up���Gʹ�Yη�u�漓�����1�w�UlFn�@}��>�P���ؿ1�ư�Z��e�ݓ�����7S�M[��U)2#Ȇfb��@?iV��6e��x~wQ^fH��q�K�VKÞx�� D���a�/	-2�Z\���2��lv�/�|���e�[���$}��e���s��7�-P~sŌش6�L'�S^, !M-�����0x���ܵp�`\�����`�E�i������{��WF2��`2�:���Ԭ)�����;G 3��'W�!f�$}G��bhIi5޴���!��y.܎��oM�6�Е�P��RB=D��[�3�Jw%3�,�Λ���*��nUe��^)����9x �N��?��b�ꏾ��p\�+��E-y^�� �`9JUGb��S'n�}�K8(FZt�%��s��CX�HQ�I �X�ob���5(ru��1
��������%����﮶���7��F�}���aC?]¾8��|��)}X�/vظ���B;T?_��35���]Y_]�w�ƿk?�[��R�͆J<�Z��¹�0���-��1 ��I�Vb�֔��2�9�$�9��G���3zq�iD�8�E﹉�F�-�a�-a"=��Di?2T�c��hk��p4x�~�"P|]&�Mžƚ^�ei|D9K���ƣS�T��ɬD�4�=�Ƃ��*��Z���9ԭ�j�Ҫ��-يKn�# �uF�d{�*C�4��p��{�B�5M�p1�F�ZN����;3�U�K�sB�c�Ii5�ZdC u�G�4�JIsK�Ygk;Q4���Ji*�����Ta@Y�L�s̙����҈��U�Av�������*$=߫�}�zUBF�(��ϻ�\4����Q�Z4~R�����p�Ra3hN2E���>���OJ��<�i�~�����`�ݭ3�D�r�ivBDb���w}��=��D�m#<bQ��w.Fjo_tǊ@��O�;��QBe�Xã��f���Q_^��������+'��N����:h��%�&�U	�[f�z�Kp˳�I3�b����	B�Z�K��Ē�^��)c��H�cP�����A�h53��j�Y�J�Z  +� ��`�I&�H���`�o��
��\E�����^���8�t21;£p%J�gJ5�	��ՒN����P�GN���>^gz~�1�
���w�ū�=~��n9����WvݰB���{�s15T8�s��V�>6�m��7x!�������1�џn���p�P��s�du)�ߏ�r�	۵�m+4a^��72t0��1��ޔ�J%��&6}��r#����1���$�Pi�A�H/�b�d�jE���X��jlNYm��]���P�+��p{ޯ!�<��ޕ`mC/�Y�ͥNM���}s�a����% ����T�״v����;m�)<���7�h���H��D��ɟĠr�>46�}���P��l{�Hտa�mhj����v���,4��\�U���G���8�ŵl��j���]�V����-5�[hLƖ��,+��qײiu��̜��y�ޏY�Uɽ�G���JK�s) 8�t�:����`�� X_�
:QuEO\��V*����L�B�ծ3h���W{�B�N���j����2V���F_�w{��V]QQT��Ӓ����M��z�B� E��wg�<74�}��O�qŶ��7���-+^��g�k���(�|��v���=~��S����՛�E�N_����C=W�P�����-�qc1|�;?SH��]��j���2p=c���ݎ�I6�	���ͳ6��d�c�2�Y�QJf�:���������T�H��c�H�oǚ@���d��z�&i�>���eEAr�c|�A�W�]��%xe�ʨ���;0j�i_��^��q�j��OzS,��A-�ı㣍{�8gv.c?)lį-0��sM�.�U����5�tƽ�ί;�%���~+n!Q~V_͚��&�*H�\ydrW��B���6j��8=���� �K��M�f��>�>�R�٧i)W�-��+i\���_/9��L磈�)����P�ee�Xv?=��5U�!�E�vy��A��Qs4>I(CrA<���S�w�K�Ō<�'�+�y�A�\㒥�m��|-��߫+QFw8�"�K��S7I���̺�).SxV)��~OK�OH��_SӠ@뀼O ͅ�J;&U�	�w��)rhiU�o�~�_ځ�m��T&�[��]�)nV�e�'���J�_��2m������aS+"!��ȧ��7�������j�^�P�݄�x�p��Հ��y������0?8k�6[6��ߞ����H����*���s�ٰ�,����RA�]1��b2
3�K�ć�Ɖ�n��>�����ܕu���6� �[a#�e)�wƛH���,(��]���.GF�4@,�U"�g��MfF�2����t�S��\������:Q���8�cŠ�ؐ説)�[tN�˖3��ꌜ6�/�[����?�J�[ s�k�\�l�>ɍ`���^��Y��4y�Y6�:��p�?"�d�N����?��F�z��{���J�n��7K1h+�`fɔ����B�^��Q�@2!�;��0�p�%9
7=�.E�s5��܍�)�_��D@��z�-%��M ��������	%���~����l�r�CE�fP�X�J�3�F�'C��x�q�)i=z�d�j��aE�������v���"\4�˂�[��3ҧe�#�6�������£���t����U�D�0���x���V^	�E��h���GC�1�CB#�xs4�\��a�T#�#{p�H��_B�	|�%�4L�;� a�
:�R��4ӆ~]8 �">p���>pa<>rN���4�N����)��(��
~έA�Ҷ�vF��y,*�_z�#9��j=i�n�;���hN�˗�o6A#9-!��㜾xK<���H��ѿzZ�r2Hm  �Bt־��A���E�|/w6l�r��c�۔�1�h-H���s���&<殞W���bu:�i�fB����.'�g��F��q�Uga1���-&;��=];�-!����L�_r�[0�C檦�T�HP��Jӟ��!'U�U&���Yd�+u�'<¾2�^?�?�n[l	RM^э����#�(������|j��s�}&vR$�����p�Gt��gv�������<��U��"�q� l�m׫SH��C�ԕy��j�qC�6-�1e��L�#�E,��3��J��m-W��X���Q�x��9{��/F�V�{M)����cs`����j�'[3a�(��,Q���Fxq��՗�zN��ƅ���7)%��_�v���J�i�ߞ�qt���-�1��3�QN����n��sF]����?M��Q}�>�p�-��>x�S[8�^�kנ!S��|�e����E4R}O/&��MNi�]�B��hpn4��C�!��=ls�m<@^���y�SͲRm��4�i���v�c��h�C;������%-��=zېṔ���8S-�4�`/O��8y*"��(�J�.�PqZ�MT��_�.��߃Rp~�>j��XT�e	�0��g�LNi��H��A�C&�|�f�c㊉���/�ɜ~���d@�	��D	E��d�<q�t��s9l�<������z��{�a������.�1����,s�IA�0`�|S%� 1�ݔ��G�sH{��J�Sz�[y��@Ѱ�޺��{�@��[�C�r
̈��L����g'�Hf���h9[Q[Μ���R����Vp��Qz�{�5�c�Hm�<�H��/Ye�2~�����x�EeB_Frɱx\��.�+�� vB�� ��o�oD<�-�n6��r��@��Y��A��+�b�o�	b�^U�/]Cfhm�i���8#J�k�fDc����c��E�wM6�W���}���Urvc=����\(1��c �~$\�x��F/�NUD�� Eq�S߲���#6�[��[h?�*��F���#��״�і_H�IuC�ѿG�n��܄4��l���?w6��ڶn�	�c��u�kD�v�cJF������ʤ�qā�5su��.��h��4�o����uP�$�(�iF6��$���%���9��o�0��/�9#O)P��'��ǿ+6�xEy ��ͺ�C_��1���H�E ��yF��(�ɩ�gʉb�4�Ԉ}
i>��0�7�.��9�2���wc����u���������<h��T�	��=9o#`�w���!�9�n�����n&w�Bƶ:g_�i�P~a~ʒ̊}x��=��0��#���1��A�H����K��-�[$�b�Z�O"�Z&�{W=�:�;:#�k����8�0���UҺ�c���gI�z��{Y����ý�yJk�|Ag��k>��GD���&�5�3��qt7�I j�_-t�#����fM��a�,��8_aՃ.�#3�����n��T�`b�ÅpD����Si |��`]#��AZ.&pZ{���uO}X��k��f=��K�QL�eؓ{��gL��-F����n�H�w�\�hdt5�E:p�v1�U��{XHyc��Xǫ��!H�ٶ kzgm����؏cT?(p����d�G�PJ��W�I?�����9�;@�{S�|���7O�-��Ȯa��6T�ﶽT��G&a:߃�k1w�(p��qiiqmqw*@\�:��w�����EhN8�?�����86V��? MQ����2T��Q��H�L7n^y���rsY��i�q��.�]�+�}*J���t�r�X}uȇkPpef��0�Z=�=�j<,��=)���]�ٓ̢"���9��S�5=��k����k�=�3a5JՅ~�,�חR��܁����U��%&�����J�?�[alq��ʑԯ���$��t�)�A�4�s�=%�z[���=*9g���߂��~���(�����{��Z���s���(#��s&���ـK}&45M��D
3��=��i/RQF�}E��W������|ͫz�g�G�����h��^�n��NŤKK�jN�/p�S���DzHj�m���0�/(��En�������?�(U/8`���uK��q�JMDXp��x톇����>���w��[�Q�G/�� r!M���0�u�VS��^����.�x�f�6�j!��&u�mD��'���@���5��jɰ�X"bJ�^�5i���N\ھ�@������#'�K�Xu	��D�@>Kq���e*��9T.*�h�F�m#Bs�����g�1�?uE�)�_���ׂ�����_1��Е�](��<Xɑ��Urږ7�!6��߭K�s���۳x6�%,��	�H¸�(��in�����G�!z�N�j�u(qc�p�ha[�v���ྌ����5��`� d�1�Z���������|ȭ��r���ع���g��#JƚB�kS�M	B�Y��`_Bգ�/Ic�sd�Yu�Ȟ��5�8<F!P��`>����,�Q\�X�5��T�{J/v�t���$Q�/n
�c8^��g��/#�(��X[`x,��lF����ґr,s =:�q� 'g{*��M4�Jm��I8�&�A�v���.��_<����8c�|���Q?5�O�ڋ�4�����؟P)���^#c'���"���M��|�$-#E���'�Ȩ)+�^>n4����G
�X�����OC}��L�s��#�VL�>˹��hv\�qɘxؤ4��^�DV���'��Ӊ�u�>��S��_Z����'��-{��\�dGE�H��L;�Čb�>ʩ#PU��Q�9s��k�0�~���gyj�>{�X����!p��`��{��}LF��zs�]� �~�Tk�P��>�]\��8Ǉٗm�$��E�49r=�������e�z_/m��72�j��	<��A"�5�D��_�R3�(;���}{c`	8��N����.��A~�:���ƀ8D���e�S��T��������-���d2	Vц��x����dm?1���y	�#��!Ҕs���=t�+y����"r���H�?�Q�?�y@ὴ#39�:�W#Cuh �{��!��m�c}��k=��-z0P�D����ƄAM�_i�C���ј��:��4�. ��[~cOo��O�gX��g�<�?Th㜩O�ϏY��7�\Ad^��t�|
����('D��b����U��싎;1��e)�ds�����:�
:a�<��J�=�����'f	�h��FN��ׯЅ���#'�bi��.�Q�|C��c���s-/di��^���egܔ-%�؝O9՝{t��5ƾ�{�n�V�d\�Z�!I+��e�u��g��pn�G�̌y�A�qc�7��I�<�k;|s_
5���D�%�LJ��swM����3N��+ME1���cO���(�]���Z�ZM�"�H���]��M��C��=VJ�ꩼa��4�4EXWg�|�	biZ��i�C��q^i�融��9�|5B4�/Ey��XM���y���	߂�R?�,�����W�*Swl}ؕ���������|�Y�H
��m.��[����3�zR,�~��T�w�
�]�i0@�BS�8+.Z��k	C�x������|x����Vg#t�mP^Ͻ��^���/1�/�л��
3߃�tt^�����ʢ*��o=+��4Ё�����v6��~C ׄئ�{LP}����Mf,�B��_��u�Eguv�b�e���C*���s\s�dtUC���e���Mvw�4o�j�Z�g��!�L�)��P����z����
fj�Ήw�	b�X��[wK��Zg$T/��Xk����ݒ�	]=�!���*�y�R<5	���R��n����mj��%Ԛ���-}��ك0c�A��Y�}L'�Ȭ�X��?���<o��Rh7v�S���G���fG��A@�[���0#��!Ǘ�U�@87&9Q?��YO�";�v�Yj�`�ql�66j��$�8� o�ҴY��^�V��O%Lz���S�z�u�)bbq<\�9�x�ܙ�G�� nr&��C�9�aw�2�V�z���Ӹ�/�?�e��]�|�&���o���P�0%�X�����A�zg���w�i�u�tv%����ʫQ��o�� ǀQ��/x�!�}\^�L?�dݨ��b�	Z�$��&&O����KoL�N��� ��4q%��%�|%���z�
��b�� ����u� v��4Xc�|j5�#�<���tN�� �+�%�P%�ߡftvP����Y��7e�n��c?�=m������:�4�aDU�~�3v<�lh,�!+4GC��7N
��DYZ��I�Av�5[������MTz��L�l���N�:R��M�g!�.���_�"A�C��^�&e �TiǓ��ݿLf�bߙm��J���/;Xx��R|ۃW�_P�S��+�k�q!��%I�Ii� �Ttn�]�W��:߭Q���X���^�ﲄe������%N�k���4�?`7x���Ꙓш�'x]y*�o)�q��ҷ��.mD��_U�$)N�h��1g�>��+�u�e��bF���-���`<f3�A��17�A��"7�8�6M9�{�&<��@�=\�������ܩ��l�����os'9�d���X'&�oT���r
����."<s��4]��:%���k]����<��'DK>T��Dk�1]���N�|��<]�ǘ��~�C8�
�y�8��mc��B;%"L8��7ܸ�[d�e[�>���?S����4d��;��v�53�'����b�q��(��j��;�����1��w�B���_�R}N+���!}\��	��%�^�;���L�;��ru�kA����.&�ث���/�1�/Wqt��iC:��"�|��H��4�^�_�Ͽ���LKe	�;�[�lu-!���E�S	u$̑����~T&�a��5:����_?��If�q�������yc��/��U?B�z���;�peIV�e�#B@<|&Zs�a��	"���)���8:���{�nծ�0AMT�X�	좍�G�@�Fv���D5y#��g{� �)��K��YMVE�G��s�Qm>O��r{�O� �]��"K��JA�:h�/��ٴ!.qE��s#<��*��*�r���0�U�a
"�&�E4�(N�����ú�w�X�����hcfP7��ޮ����!� r��'T_Gw�"5 ���hާ�,w���i{�0[�Y���!ˬ��u����ä�/����}�������O���
+�ʑ.�zO8x0��C5�,�W=�+5���셓؆$&[��K�� ��e>�ny���ܹZ+&�u_+ap�� �]	�G��aiaɇ��.�k�Qn�UGW����T;��(`�������lٛF&�E�(u�(�Hk��	&��^��	��P�a��>��$��k����z��כ�:���H����@���6Y)��e�ڎ��}Ƃ�ɧ����} ;�V�f�I
��C�bU>�D�^�s8�$#��mI^2j�~;3%d�ë��k��3~O6��C.bL�� A��"��y�<�j��`�O��������AgQ.^˶]Y
�3�z���iK�Lf�4���Ҷ{�K��"���@�s(6ë<�
O��3#"]��}��.���Mq��� S*-���ܦQu�n�J^�L�=������C1L�
s[��Z#kM����t��kQ(������}x�a������~�w�F����x�T;Z�2�J|I`X�R2%W\|�j���,ׁ���d�V��I^�%8�@P�J�ҧ/���UO��'�*�O��;���p�)����j��o����S�Ո^1�,~D4Po�)�H2�w��s��ӈ��`�#ѳ������Vp4J��!��J.Q����ow��Tx��'�j�H�j�:�[g�ы�NjTB.(l�����b�m#J<�T�ς� �1>�T��}��b�;E�C�&��}ȳ<a��Ϙe
�HW
׊��Haf��U�>���u�S��b���`m���|+E�Qq �9��.yrA����֤8��O�K A��7l��4��F-���y 	�\��CDr�"
Rd��Y鶅ũ�f�,�d��n�3��=.�u�l
b�����1�F��%)��r1��jm	&7X�����(ލP�\h����,Sz�n��\�I郊J�L���zժ��>��@�f{��8g<<!Q� ����b��<4W߀��dJ�8���7�R;·�PJ��C����
�k�y(�֭~I�eϨi8��~)�x�) ���#dEE��m�6Z��)d��ƞ�b�+�j+zTwM�hl�m[ F@&=Rz&�z���*Zv����&�=��KxJ�	tʏ˥�}����I5ȶ�{7~4�M��y2O�7)��Q/٩K��Ekk+�V��m>�ni��:{��H�|�o?&~�'굚d�`�������<t���8�2[�]�̕�d�q����
�/������= �&�AUzGu�Woʓp=ULҌ��Uz�z�#W����=ckww�჻Pp�R���H+�3�b�t�&T�^��ծ��Pf���X95��8u�ҴbvJt���:n����I���9 >��J`D�|BnD{�]�ܴA%]���Zl�Aq���I���8�6��b8k����P	#�R(�
AM�MlGꅝ��H�9�4������MQ���Ň�X40s���x����0��H�y�?QC �/��r�
����ᙐ�`�k�$�& ��V���F��qLt���g���ـg��tt{�yL݆	��,+��8a���S����2QM�5� ec\t�.�Qw��@Fv4���%���DA����'�"'��կ� d�n�7P��f�q�ω��Z���A9���.�/��[vW����]�*yG q��=���^W1�Z���C�\ �m@�����]��w&�[v��h������R���|Z`�jE�ڗ��y d��OCu@���Jᲅ��0l;k�U��
���wp�`�������&�qԶ��;;�b�f��:t�:Y��Ri.M~R�\��nE-P��<aw4]\)jF9LNLp5W��C���- �ˢE��y�V
�.Z|a����HRV��T�>s����ӟ�em��'�*���^�HZ�]���� '��
�O��F	��V��3��֬Ar<qv`� ���$��d2�`�$}�v.�v���VT�>�:�h��|4��yO?h�D�9Q �aqR�wN�ߡ������$�Bw ��!��6�K�$膎Z���Z�ޡLk���[m���7�(խK�+QУ]��#C�\�Y��]����X��x�7�]���:�I�H�s�FQ̉�|o"K�ˢ	9�v�j��W��[~�V��cp��`��^y9=������2���s�E?L�	M����0�� �BZw��$�56s*� ^l�����7נ�J�D}����-i��*��O㹪l6�|��_�����|�N^����k�g��_�M�����S�'R��1(�-���q��i=4��m�(NV	l���p�j�HJ)l�Hz�퓫�$���wJ��i�E>�j�P��o4M����֌�ad�W�\K9��8��AC+��]Nٛ����� ����n�L���s�^g�)��V(�ȿ��v�TV>�c��*R�}��ܟ�BNY�e����'�i����uBL��I��X´"�SP�µ(���<Uc�'�%ᇁ^g�䳯����<4.p?������ ������N4oGG������\��,�j޲>�'���Wl����.�����W�I����a�� �P~y*Kދ\�`}�9���P����Fɗ����Z�Cb~g)ֿ���\�:W����t<dt�����Z�\7��QK&ʥ+B�����f�=H��\P����.�Ť7�V�	���L4����P��?6�����b��w��}Ų�8Kɲ�����u�0t*�����l���́�O?��/�l�Ns_���AQ�K𠫏��gK����=Θ�}Vq	�hQ^P��V�^	R��,��VV�^�C�`:-B�S��=���Ϝ5+3=����L���r�U���/�4z�SGR����G��������8Gdh�2���:$�G�X|ldj���v^!F�N�N���lս��}ݰaR��9^�����_�V�رo������[� ��+E����i�2�����]�Ĕ5F���3S��x}61�����Q$/��a	��_YT̩�L��8��^61R��T�LM��4�-��kДkw{�d���?i����ߙ���劒�HnU�	�R:�@���v�nu6G=Nā�J�-@t��)'��i˸Q6"��Fl��^�5<�-�T�O�J?<X���ua�1���#JN@��e���>*7-�����	["nmX)X�^�9�o�2�)]���6�|1x���d$�fOql�|&��X���b��H��)m����"�R��Hs���y��LwX��vA%s�1/f-\��N�����6Ǟ���ap�2�� ��ʫㅞ"d	.�xH��w?؎��9�r��nڄL1Q�'�{�b�Ok��K �]��H���k��Yܦ!�:V�W��Q��,!�*3�`c{P�w$����L0�m�r+z�F���=��ӊ��G�1\����)����ne�iy�&r%@�f�ƚ+��
�+���eH��@4�+CN�z�&v���8�D�J��?�	�x_��1N��t�.�% ���^YdL�tQI�!`RM���ii+�CT�o>�z��v�+�\v����N���:�R�F��m�
���o���ōXQ������ ��ӐЗ�~8�@�qR��	�CB�z
|�nU��.�@��2����.H'1`%Yy���Ƶ���^�u���}oa�^�C19	�*��qz�g�-dziw��F�ݙ'�-d����"~'sS.��۶jK��+�I����b��w<�]~�jJ�½�נ���Ž�M�s�Lc�J�K/��������|����Pq�ue��|��C/�� {�����Sq�-�����W�E���$�~m;�"��떓ñM��~|�)L��.�7c�5��.���Zz`(�����7
@��;G)5#��E�q�E����Jn���-�$�>���.V�J3oT��|��,��Qp�$�7���	��7�q�����-�\�%:�_Uǩ��_=h�F��+S�I<~����(�L���E��|�vR�ﯜ�~�e�>ջ{��-9EV%�1��&�	e���8�zz���_bL�юZ�t�X�ڂ���v�U���ԦT����Az�E�J��N]��Z�ۅ��\Μ�!罬���c�i"��Ɋ\"��f|}�32�z	��[T�gc�&�ȱ��'	��9W��B�^ΞP�r3���H"�&�"j�̠�,��!��h�f?�G��������!Ѩ���\����?I��Md=�D��؅�=>�W�ٳ`D��N'�HmL:�V (h+C�:*�s����H�.�I��`�Ϯ =G�܅���z�>��L�˽E(O���#<ȏ"]b/B931�kДi�yU"���w����u�1'�E�&&�~\Cjt�/.Z0ۅ�C#�иT��:�!d9���-��K��$f>-���B�"NתN��0�˙7 �.Я����X/(�"�u�f�sJKpI3dj��_��0T�_w�z��d����g��i��8?�/ޥ�+�B~T����3�!6��*C���d^9�=�Tw���lQ_t��r�<z�\.�2.{I��C�����qEg1�B����:$����p]S���SJ��vL��(-�p�&]�su�7�[�0>.��IBa�s(=��7�[��Ō��x��K|7)�o���|��t����T�_��ؾ�Ƚ��%�zGW	#7���J̥�}Q�*g��3���g`9~�x@�Y5�����[�sta����t��/l�*��Մ�ݪ�,�C�ϸ���@Y��F�x��-'U�f=n)���*?�<��2]�^@���Q*e��1
�+U��nV�����Kʍ�\Ry���P�l���GOy6m��&��'�)^�����L�p�����U�P�<��oi�c�St�.�Q>��	�R���L�Z�g�r-�6	5�8�I|"�.�|"���?YX�&0{���oOEk�5D��B���Z�0�f��ĥJ�ic�w���	��q�;�a4����8��Ό�:�Z8�&j�)ڴϽg.��HJ�_��VO���P߯78��,��pL},t8<Ű����d��W�r�HD��D��F1�l�4��{I�.�Z>$[�q�{�7�_��g�Q��u������K�N���Ln�4;B�@J)��ǒ��G�u]J�B=�F�,&gU������k�M�Ҭd��V��+
-�l2�)�;���oE��X�8|�d���]�C����dbN��W&{�؁����H�w�;�Z��C܆Ε�ݷ�#Q�6b{������WZ!����d�����]D����� ���3��O��/���9��.�"�U��yO%����5�e�̠GU�L5T��D.Е����O���L��b�O���J���r
�\:r�_eS@DLV��8�6֜+eya1vp�ih��.x?*�p�-�����pKӲ�Tg��F6�D��|�a��Ĉ�#aJ����6(�-��J���e,��+5��n����9Oj!ba�^�F�����Mv.��`��DD�d��M_�5E�����v�����K3I
ZAG�s�IºE�|z޼�z#=H ��-��qk�*~\o4~Ԩ�,���횤�s5`�Ժ+��&�����NZPތ�ti%����#Rč�/iӗ�-��!�`�O�o�I�jRl���|��#����Fz2����o`����%�6�g���=��x�Qɫ���*�c��ڗ���j�"F���0(Y��U9 ��*����{F���{R��_�֠�+��,7Y�Ր��W��+ܐ[��k�7$����5��}HV�<g�/�i�X.�᡾T�X�������)"Q�Í��{��d���0���6��y'8YiǕ�&,�ժ1!�Awc����� *1�Y��i���ة;8�ku=F�L�� ��t��w��*g�����/t�Ewy�Ʌ�R�#�`�'+2F�Eӡ�ШEbT�\]����{Uޥ���fe8(�Dn��$~n]%ݱ뇥�5�5/uԢ+�����	f qc��L�_*2#�#8�-��%��<�T��v�`�yY'aF���b�=�b����+�0�e1��d�I���
�k'�Dܶ=���=³L1�M��H�����ǫ?P��p�",�3�������R�H��|rN��]|��5NI2v�.���k���E3��Z�5���	���O��þ��[��&�ӝ��ɗQ.��������=�Rvl� ���ִ�4<�.o,A�����U��O�p�pָ��7�p�lM�z7�T�G^��3暈_��t��w)��BrΓa�~�+���rD_E�R|��f� 5�1Q��<�� ��)$��w��#�� �W]:Z�[,�<b��H�P+�^�+���f�b\|���A�T������bm�l��	b �MB���۬^!������Ƴ�`Ā���Z�PT��՗٫��J�;�։\�X^�"u(�EO��}����T��4��s�;�l��ap�n8V@��TՔ�����:�ԩI�kp�����s��f0�J�=���-ݰ"K�F�H���23�e; M�?�Me��Q��G��,n:�o������`X��+AR���(=&�i��=���*D\@���Bة��?�������W�;�3�G3ں�[0�#cn�,<���9���l����M[�3����B��gw]�������?����x8ez��l��w�	v��uRBM�rw^ҜTF��0ƕzvsb��tRc��l_���HhW
�Ȁa�y%��}z���+��z�Y0���ʿ;��4���͵��"V�OeÞQ���U$��cɵs���_�/�&%C�@f'����nu�:�x¢/ɢ���� ˰ �
x2h��*ퟲDE�I�/4zz���j���m�2����.�(o���S�:��?���?aul�������� �HURw�C�R�ņ ��R�e�k�g�@J_x���M�@�L��\�}!�gF�"��xM�
ڤ����֛� �̉���]�j�2qM:���]�/�WT�%��9d��HG[�fӹ�S�EYϠ!�����5̻�!ݘp;�t�3�/ݠ�1�9cR��,Rhų<t�9���f=�e1/=�\sy{�jD���Y���[W���y��e�&=㣶جߘv��g�oH��e����1.�9T�i���ڌW��p�ܠ�-�0I��8��ʧ��v1EjM�&����Y��˫���s�B �(ݦ{;�A$����8�#ڞdqG��·2�S���0��=9�]�h"�A��)	�`:T��"��ۜ]���U�P]�p�7\p�"�b'��8����n:�e��,�F�ح�`~}��Ɵ@��?iT�CD�a�(7�26N����k��2 D������|����,����uV�t!��8y���F�rO��6�p�j���/?�+�'hǕl�ς���f�I��Th�uFM�Y�������a���[����'D�pǁ$�g(	SF�P�Å�]��U�m���M��&���Y(C�d������V�@T}f�-+?�AL�V;�n�Ea�B��E�{��*�M1k��Il$���MѳU�M]"�+4�g\�K��ǖ���l��K��RR�9_��͓�p1,n��s{zYh�V}��H���i;����h�Ctm9��x�b��1@lW
�-��L��� ��:>�]����LŢ�=��M�I�����W�����<>�f5�l\�G���u���e�_�=���f~�������D��IN{���~A{��8R+��hr����|Q\u�*^ ���_���9@"Q^a*c��sNY��c���*AS��<N�"L��I�w�}�mb������ʯ�MC�-�w���V�B�V���!�	Ц�	�P~&�c��|��yq�RFd��г���>I�K���-�,jWL��>s|���HL{�'\�OAa�� �]BK��ࢱ���37Z#Z|F�o�������[j�	9T�[�ށg���VJ%�tY;rm��h���e05��0���F��I%��UjR����/(���d��
]r�W���H�}�;��Y�5���'�h3 O4�QjZޑ�h�'��.
ڋ�kQǮ|p��o�fS�x�ΫԴ���a����'�G�>�P�i[*��W<���,���/.[�@H.#�RQ^���N��(.�2�m�P�dHO�)��P���M(�!c�13{���+ȅ#��3���� ���Q&'��`H[s5�XEE�4UK�;�9��cWذ�(��h�.��� {��	6q~脈9:x�y�����es��_��|]�3΁�|DB��hr��^e൛^�B�e�F  ˮ�����;�խRӁ�E�g���G�u���D)��`D���L'z7�v���>�b��S�s�7����<��y$�C|Q���}s�h���4B/ź��yBf��z��ϮΉ��XO;KŜDvN�N7�=Ǿ���/�M����K�n�k�Òר��):9@R=k�ҹ���3�.����Ġ��Kә�6���c�� 7�'}�~;*�������%�}�-\4����^�]�Xs�Q|.�ڬ���!t��Dft�ɛdō�\J�yM)�4�ߌ;�����[��~iC�<�&�[2q˗�PmW����z��B�W�[����v���R�<P:!�1�E�t{��uB����p/���%.=ªZɀd~�(��r�bmk�۷>\�����V��\D�׮Y��	�@�]� ��h���e�P����
I�/R��Ci
�~z�~�yu;����C��-V,]l�4K��	8H3ߞ��*&������5��#c(��2Yn��9f�f�3���ϯ�W���!Q�u�B�yq��X��z�!ul}�}Kþ��x o�0��P�^�5�,�AXW�f�1��u�g�/�#쬜,�FyGq���f���c�ot��� =�� ������_�ń�G�������R8�j��e{l1�[u��%�4�~9=����c��j���ǧZC����'1*�^-��]05K�ٚ��I���ڋ��9o���$�3B�=(���a;0B?��)����~�����D�)BJ"ζ�Q��
��M�l�4�o�Sċ����s>	!�ŘT�%WUr�P�̷EËB�$LXk!����٬��'cU��Ő�J��~��|���]��� �G�E�ZH+�ve#��aM�3�jH���4�Xtx�	�)�іL�4&��L#�#��y����)ɨv���Q�tj9&�g.vcx�*�İ@T��T�F�]o>�u�"�7��s�X�ۦ�/���e	1 �2KB��p\���������B1 q�K!�/�6R���T��g0�?�����xK��)�T�f{�0=��Y��gN\Q�\�Df�v4���Y��&��I
.#X;	Ux�?��;kԲ/��^�31�����X��b����}�H�*�U>���&�B�������������Bۻ��8�*G�zPJGO���1fY�]ێ��F����}m��ā�\|�Don!�{��X�
������Tܫg��MR�?�b�|��+���^N�E��b��Z���W��׭����珽Q`=$�m����ܥbIF���{(b����z��x9��̣��$j���G�X�D>�h'�׿���1���c*����;�A;�C���ᙕp.7�4V�I4���}ɲ1��Ե�U6M�;
3�8����^JE�q!��C��Y�r����b��Jxy=�\�0%�2�J ����D,�7��f�׫
C:B���/�Z�՘;���?#;��u�MS�(��u��c�3 p�s>E],<�I����ԫ"8 e�SUMx�\�DF\9ێ���ߝ�V�L�w>0S�`T҆B��D9��X��[\������^�4Ib_�+f)��^�^��l��_�$Utw�K8�@=�[\Mm���ǲ�=�cSt�B����� �{Q}،�8hj^�m;A�o9$�yH�V�wƎ!�$���2���8>)�N�t�����^�78/�2-�qn�]�`�@�Nc*iP䇟�4�1_��^�5�RP�)�#o��e��%W�Ƀ7�CڥA�˜MHFd���'�0��I�-A����ogX(��qj���k�=~�b��=W7�M
����F��h���{6��*�Te}:/�h"�<Ԗ8��LOk�;)+�RN�i��r��o(����&���GrV��)k�� 7]��8{���l�-�j����ZY(,�7�V�r2�#_pWF��|�8r�:9D���"D	�tp	�|?ki\ø\Q�&�����4/����f�p�Ģϳ]M�ú�T{;�"�#j��\��\<�� �&g	�E�v�2k���r���۞�j��J�h�C4տ� ��ή��x_�n�8h�6�1�|Yt]�>��V��w�1|!c�����|�gj�����hZ_w��Ng�э<��U��A�#�R�����w�o�T��	�th+�b�Z�̤A*!ų��8�~�
�F%\��b�Ԗ�7"?�_�&wN�Q"	�T�~��F�Ъ�!$�z��nXI��ْ��/�b��镬�XiI
��uR`��뉷-?tz��I�����[D-04��E��݁r�c`&�z>h���?�j=�������BR���FW���N��v�y�?2q�m�;t��#t��pwTu��R�b�㓆��b�M������=��ڔճ���ϗ��p�9�d�Sr`2��Ȃ;�}%_{EҴ��
5��ڄ�=<0������0�A���rE����!���J��C:9�I���4i����u�����0�Sl%#@��<Im:��5�i_�ܬZ2�/������n�$�]7�'!N� S��qA��^�.R���*��C3��~�[�g��@������:��+S�On����Gi�3o�d��W ����Kc��!�]�+��h��B)�ц}+�H&-VD!CzM�p�t��O�XB����l:�?\�V*�_+;}��7��p���J|
2�p-�����H��0��1�h	���_���[��3��ٴ4a"ʽ�����o��f��Dh�61~"6inQ&5h����B��p�g���5٩��8����Ex"'V����7������	6x��vI�K��b�����D2(��5/��'��_ )�U�پ�ApM�3Z�8�A�MVs.)|��>T��Y-��^�	/?��{�%��s"5C�[�\�4�6�3����4ҫpSd>�H���a#ߦ�W�%����MWJ��I�A�ȱ�#q�D��.� '�+��7�)U���-���1��ʹ�B��/��Z'���з��-���95w�ᎎ�riVZK��ү<��>���lr��x4��|Bc+=�>���h��}	̄xS�-�ގ{�	��T��gm�U7�9���J �]ǚ�,r%6U��5`�.ۮƏY�<|�����۱2��@)l�ꁕE�bh %7dr�I�ڢuh������  CZ��KgaS[C7�7�Y�<B~IDF����͆��mv��Y3�kL~x�3�V (���)�5��{[#Qܖ�55�p��'�Eq�nB1�Jo�!�Y��%��xEw�$��_�#4 ��C��H5��$�9�h0c6�H�F�R;Wp"n����&���uW�,�3��L_Gǌ2�#0�C�c��ʓ��Mޢ���vPj�ֵ�A�A)�ˉ��~ie��+���q��n(���'�\p�&@��rc���&e���[�&B	�į9������b�<<Ja0��B�C���u�! E*"�d�w	qN�sѥ[<U��u��d ��>��|�m.f��l���#U*z<X�E �v�ե��B���ʐ�9&z��ut��_s�r�w���j�<�[G3�kE��W��m�_V��|g?���w`���@�bs7�����e�N_��떙i
�?'2`�}Be#t�g>k
]xw=�^��X=��S|�H�|%}ө[�wS=�-���sa吠\KoR��)�(��iO9%0��8K�ļ*!��Oi��7�K�����Z�� ��#,��7��煓]���֦��!�i���]{����)�l?��� al�~�7��("(�f:*�	x� ۆ�p�a��gevL'��J�jsA_H^=��ڳK�~��Oa)���"�k��Q/��Q��λ˦��C'm_���<&K�����t�|m�k������|.�A�õ,u����H)�&ⷡ�V
�srZ�fؽJ���W��_04�PT�Pќ�#����x�ԠNk���F�OL.w�"��SFD��Q��z'�P��̣Ӫ��(]W	ބ(���At�8�����1B�tC����d�b�%�Y;���ӟ���%GjN�`�Q :�3&]�rw����P�K!�-�!>�Ts�l����Q!��V t�?R�O�*�NG)\;�:�1]V��k�c~����:��}n(�e�����<mp�Ӣe�`�?�؄��OD܋D]R��I�s����Hp\�F�ȱ6ˣ�c�][,Z��� U�#���}LFp��Cf|��#�7)�D����i��OQdqW� e������������@��֝�P�>"K��!j�vۘ��{:��>��O/k��&�ɾ�#��{�w���S��K�9�%3Y��1Y���9�.�?R�m|T*�c[E/ʾ�+��=m�,��*���\,�n7�AY���ohRIo�:���Ԩ�W����_BmM�Y@�Anfo���_�˅Z	�?'N6i*ŊO��G��eS�X2���AT�&�yJ��:΀jZ%,m��(1/Q=4�o̥C81w(Up��0��d/��M�S��դ+�va��� ��ģ%�1.�)�
I��p� ����-[f��C.`Ȱ�H��߄��O�}���V��Ɗ�f���|�&�Q��1�\�4+Z���}����&�)�E\5Ȑ���59T8oG��H5�*�K�QO��8�%���{s$(�<�"O�b�:������Yj���D�(�F.�K�i�ĴX�ut&ȑ "�ع�08����{��tAN���QT��!��7�\)đM.������c/9Lu�k�)��� 4�a����!���/R�k�V̑=�$bܰ���?�,a��HL]x��"f���{�3������Gi���J���W��N�RgXh ;�3{q��H=a���>�.&9�����M�2���k7���(�Q\Q����B�t���`W����7IQ�ֲwzd�C��!�sc�2%��]���f�P"�%��\؊CD���"[��:;i�������R:ߥu�'�O�p�^
\�����f�⸬7�)ˏϲ-�}��u��	ҟt�	G�waԋ�{ 7�F{k~���h�8�]�VO��l4P`B!��6h�+�s!�ډ�9qK�[W��K�Z�y��646$Y�(�`�w���t|/��]�z�xn-ja��P��Яl¬���w�#�7]̋5h�����[��-Ҩ��F;�Kkx����6.e�����$�7��b?�!tv���h:���2?b@\�o����/6�2U�����f�Qk�w���Cb?[�g��c�m>�PrR-K��>,�&MC����v�F�'
�Dg�K5���M���G�^��>"�)XRQ�ծ�EUŒ>�87��y ��\V�x@��Q2��۰���]dE8���M�N��Qp�q퀾��m�D�I�+�U�/��PW	�Dk�)��j�v~���jj\��ߎ6���he�V�#� 1�n�>l�Uʦm��6k��؁32x v�馠�zL*��(�m] ������&��HpU���O4��&ds��tb�*eGd�%�OmE'r �ZMx�%�!��!�9!6�4����/� �9 K�9�Z<�!�)�ϟU�8WY��yc\��&�^l�-U���U��}2)���*����O�zr�}�
j�yG������9Igi����ґ���<���:��ve��?�K����e�L�@�R�����b��gDy�ע�b��#�������Ԯ��"���'�O�]���F@vn)+k" .F��+��(Xv�|ר����rr?��kk6˿EKs���z�wi�C��"R��X?�Qx�/�G�B�aj�8z�y��\�M�Ȱ�9�,�0G~��:�:��C��u��꟟t�k��.�%Vľ,��س��:ڹ��O�H�I5�1`!�����8�S((	�=��W�m-����䩂�0�d�&W=��V�	���p������D��OL~B~��Y6�(/F����Z�f+ b��u� P>�~�	g�*Y��ו��A�z!ܧMI+�QIu���aAaA�G�\�z�>Cݤ�wSry��t���x���'����5u��+%Byo���1֐�,��W�b���M~�t�����a��I� }S��G�)?q�F漉*V��6���.p�wl�c�O�
�����CQջ��)���u7P��[�]���Du�fb��L{ڭP�H��:��tEg�U^db�	gٝ�����@tL�p�%
�P9�)w���+o��:�>��eps�p�:`�O�:�~�����Kf�Tw���9��Y6X��X�?@ר-#X�D7T�������-����e����Ezk4k�Nb󞣋��>"�1�����	E�.�-9BM�,����C@��3���\|`>Wӄ:_���S�G�2���p��`��n�����X]"Do68�I��;�������䬗4�{����L�g�vM�.������	��w$9��C���E�f_.!/�ww>"��u!K�%
�,��4G�p�. 1��/�8h�9�j3��ij�����;�}�1�ɢ��Y�ko�0�j7<�K	�(!=��x�v�t;��md��d�&֞��Q8V(3E�����6	��&���3"x��4x$@%��Q�:kq�2�^;���lWYb��o���Ue�27?����(z�;i�ɀ"�%?B�yh��˟k�I��w\2��[��ME�0��Q4*6�/� �p�7��#!��1�s����Wa�)�ಶ�7��A!�D� ���賙��~q��T��џ3������ׁ�-Ɋڪ��r�n�x��֚��B��_�͇?x~g����.��'w�u��'|�肱��4���1ۃKGkeI�
��A!���97t1��y�Hdv`��{V<�uks��-� �Z��4�Sw�t<��.��+� ��nCp��bAZ��"�����f��sŠ�*_�h�z	ֵ�`��OŐϖ��el¶A����)�s�5�=�����L&Hah4�=��&B)�ş/Y�ؿ���.�����
���g\J��:�3�"��6.�^�Ķ(�ح�i���d#G6N��,n�����+9?뫱{�I��B�$(�Z�����}�.Vo�]������LCo4�1*Ǌ ^��pƝ�>����`J�K���'�L,Y&K�)�P���9�L��:'�憻��t�;z#땆M	f�N�p ��x�hS&ϧ3�N���R���g�.R$6P�g�od�ńoJ�C5kwm�+{�;_�,�����م*��z��x��9��F�2�S��cHJ�.ҵFUk���st���z��$��P�doa��0z��(��~�HͰ�f�e���JX��j�DDdP��r�;�iI���s��j��2=��T5]���0��i5�ۈ����#E�:�u�nw��؉�I�_`?�nc���I�ҤI�����"͠YBNX�{�8gJR[@@�'�i�&~��G�6f9���vJ�`%VN�ʱ(T��N�gn���s�s�4g�K�ف�����K%���C�h)����(h������$�����Z��w�����D��@z�:+v���:ċ�FK#b ��e5�����12�i��W?����˫�!o}��$��Bt���n|WΣ��wO3�Ơ�[Q�Y�%���]��1�jN�r�/���s�i�9��-��-o�a�0T��iࣰx�	z[|��B/��ч-��M�Z[u.#sxhZ��P�P�z�9�M��,��f� �3�|�Q���N��?{�6��󿙡28�n���^�`� �z��6��(�sMi@J�o�%��4j�[=D��l�ݞ�1.,"@Y�5@M��O��T@V��ą�]�}��Ѷ����U������;(
�}�Ms�p?@]���n��HF�Q"��X��cx��Z�Eωʴe��U#ϑF�H����F�u��Zl���U,�AO�WX�2���%����܅�h�(R���;�Ҽ'���u"����������).���Fɮ�A���
)0�vÿ��F^rN�ϣ���}��\2�7�"��*Y[��q�a��8�Z��&��]G�`�i���>X�H	����}ɬ\�%�=�����gG-�-%��B\����*s?���`C�Y��#`����(��Sos�����j���j:�Q$O�Z{��/&N���K���-:�z��P�ޏ�~~����=�̟�$cBg���l�C�`M��2����r�s(����>)Q���j�-G�y��q�ha��!OƾE:��7�O�����'L�H���9<|��W�H�#-�.]����v�oRP#7��za�IUj4�,�!X�O���X�o��{�ۓF�۬�{�
�mV�y��>�ѧ��x_�06�iRۯ�����&w���3pm;��C	2��E��k� �7u��#P�@V�|*K]�h��J�:"TD���d��5˒��Rv?��eh0ւ69L'�O�_�v8�AlB"��~���#)�����q@$�FZ�kU�k����©A����opw�'	_y�8�{���ݙO|]��S��Wdui4El	��� ������D�x�
�?_Fç2��
�X嚏ܱ����}��ᅙ?�X\��`��_��`�f�N}핞�I$/�iU:4tK����^8C�&`�X��pHtuo� �F"�"(�S�m��$$��-��H,�
�I���'�g�j��4od��oy�6�.��������p"=�±TI#��F�����	*�jJ�ZꞀ�ó�%���N]���	���/� {x4����)@,��1?�1�H�@��|�Q|�o���2ҝ��7��x^ײ���$]�w�J�c^Ϭc���LE�P��*��v}��zFxCǱ��s0C4?GO��l��R2	�G$���N�~z�lS�~�Ю��x��57���t��]/F�{+���p�m[ �|�n��i5]T�>�3�R��K~�+�j�_g����0*�|�y �����k�1���r���n�������.�9���a^ÜK�X�$��	pA��d�E��t�׊DyL`�U�x¯Ϝl۵(f�h��[��u�S�rF'�����KW�
�*�E��\���WE��be���=M�3|J�]�g;w��X+!n���Gq���M�!ٳษ�G���G8���{3JbP<9Z4G�5���Q��p ��v|^2`��(��l��+6!�GJ��`���v��ǁ:dw�����;L�1���8\N�Y�S�o�f��5���ī�F�euiɿz���V�4�_m���r��@Z�V�������C,�r��f$��zgA`X���Xu�=�W޸b�0������^�ׯu>9�hd
u�5A�Mr��J!YpKWk4�>�
�-�{����]{�.7��%�׵�a�5��4�V�aL���U��y}��$F�����`!ץ��t��-��j*D[o�}U( ��٘N[�we��بFυ�s�W].��W���m��y���h�世L�h�}�l�7�0�0�e޵��b�0u���f����w�鋥�ꯌ/�/�b�9\a
Z����JsY�g�b��Jw��j�=M�Is�e���Q���7.yf���^h��
͞~�HfM�O��^^��x�7������mF2�WTa�<;�Y��+6/U���������L(g���C��sT.9�j����b�[+]S`��5�_δ=��YF�tc�b��	�`2&z2�<��7�����|6-�0I��k,F"���������n��6~��ER� ���}ݪV�RQ����������kx=��9s�i�o����s��AGo�w5�|ԀX�}3]<}���@��YZv�D+8c�\o=`t��	r�Ȅ�0n��*;����)Ro����@u�t�]qB�j���s����`�+`�W	�`C=�Ţ���Zs�����'��)S��6KM��SSD����X���0�M�S��3g�J�c�3�%����ʸJnR@wʈ�x56��ܠ6�<��6>B����6�'��ʻFq�#E匮���E�P���כ6�NOp��s�-%�eխ�=<�/x�[`�&j�j�r�?$f�f��W��i@�Ӷ�u8�.�<����\�S�t�=
xr	*�K{�j)�z�������'~�R�-"`���Y���y��J�&U|� ��W�#�fׇܴ�v�T`�St�0S�[6ܓ�V��.�j�-����{�U������z��Ui�����|)�s�<��^y�F�Hr���+iu� q8V⛋� ��<9@����~�����}q�w�$	dS��G*	�G�A���:����Dj*��~
��S6��#�ԋ�v�Inl�����f��)}ꟃ�V�y�q*�=`�a�Mci�S�k��cH6��3�U���-���Xes�\�4ޗ?�:�#��CA>!C�|����7�O�F�8�UD��B��<7���z����e��f��S�7�����snv�iA�J��Α?.O(����",�6�0�n�_�n�t]�[��<T�{{���5c������i��C*���V.7��l�kf�Ԫ�_}�ڈN|,�v-7��N�"��bxW�jg��m��Z����\D�0�(����/�L�a���+��c�j��1$�
^�0	����a�����(�݁��4cq����c�H�vP�(�:�h7��7��L�g8��pst#k:�l�uC �3���p5���^Y�I�3�8��ڻ%�{֧�[��+�/�OQ�"�(O?��U�|���)酳l����%3�C��G��3�/���!q�0�uf]���7����9�C�"��J�h��K�P�BL��Α[�p�v����Om"W��j�(��6�Ũ��8�� N�h��g_y��J0�f�g'E��Fz�b5+5���>���i��7l��?v$Ξ=�R�a~\9�Un��`P#J���gH�V�,�ik9�}	�2Ǹ߯<�u�����S�&�"�|�Le�݈`���ݻ���~`y�i�����S	:=3X�������T~����ݦ�B����A��=bM���f��/Z#$*�d�-C/NQ�?���\�Q���O��f�c�#r����i�hY3fq0�O��r�B�'uj1_I�����e������*�j��-��"�����^�W0J���uE5��ɫ}�X�{����NXD�<����6����H�)N'c��j=d�M;�y��U���a�8A	<�ժ���F1id�c�,8TgUei%��9U��$.��Iu�^ft� P��m4�$q3���x�Z'�)�éBv@j�l`��o}� ��PQLe��葿�(ҝ$ss�C��B��@֖ v>���Bұ�I�z�@�,�Ȭ_,:;1=�8�@oe�%Δ8����ZD~�Y�xx[s��t
F��Z��*ԍ�$���t�ﲬ�9i�⍓���Ԍ!�%nZ쁯?�8閍3}����t5��X��B8�5�4�0 j�$z_�e*��~ :������&��i&O��"B���
��}�� ʲ�OzBS�8�և8�qN�v3��m٩{ٝMEpD��U�x�<wZSl�7��sL!�7�rA� $L_��h�.���1��Jƹ���e�M1sc.�uZ���gX$^j��*��n���£0�����l�i�{ֈA��Ni��ןH����2����m<�_ �e:N��2��_��l�ٟn򂯿�����ls��i~1��J���R����th'�oJ�bew���8p�US�
�OY�(����Z!m�I���N^ճ�F��vw��c��k;����!T?lY��[Gc��yN�Pk� :�Շ�wq����7y�V�T��3[ᱲ-�M��o��#�_���Y���8�
�H<��$������/�m8ʟ��/@p+#ִ)`*f�����U�_9��t=J�� �4�2�ԓ�/�S�D�*�ph��D.S���W/Ԡq�)��Ju�뗵jG;�~�bd{d~^����Ŕ2j�
"'�	䓈w�f��w.������?���T!Qk�,����ޔύ��Az}��_��Yԛl�iӿ�M?��N[��'ix��h�"S�h��L�V�G��&F�������{��1�� �X�[�$����;�
���
��8�OC}��!�!~����Я�-�B���~V� އ�H�Q�!�������馍�g4�&u�|#D[)!gQ籯L����	����=��ӯd��h;�W���x���M �%��O&͟��1S;��
��#ACȷf4�|�	�k
J]��e�i�Fϼ����
�������s>�(?�NI%��zomJ
�"�8�g|5)�_"���I&�k�^k	������������>��a�B�R�HPt~�"M�-p�;Es3[�	bb�o�Bh���A��2l(s�@6�5�B[�>)��듯2��I'&�:�NT�1NL�c�� ٭M���>�Sb��3��7�]����ZJ�E�E+��::�o�>w�?e�h��|��ƿ���4Ke�J��F�+Y+X�8�2�_:$���*a��<����_��6�J�wX���o�\kp�ڰ�0ʼ���8&�%���!�7�RѸ�1:���9o�j(�����{;�jm�e���m��\V�2G/�����$'��I? &���<�8�P�P��m��%YG�TKN"J%��ʝ��|�����s�$��
A��at�4��<?����!����HUi�Bxl��cBV3��'@�^��:ol�"uW䇘P�t�]P�q[¢Ł�r�~!�A�߭*�P?2%clU$�1�lV��pϋ;%5@�����$��+L�5V�:ؖ�w�މ�M�Y�{�3�dL�Xʻ��� ��m$fQ�o�Dj6�g�=�Jս������b%9cW��D?<��-� �ϩ��G_�f�u�-�����c��n.o}�rfՆ��o�Yr�[�H�'��ݿM�c�љ���'v�Uqg�ſ֝�r.Z���fJ@ݶ)F���8��O�&�=�JI�Sy�hq��#��(���=J.�E��2؄�,������� �[E+L�-&�w*�ujmaގ2�1��uʪ����\�M�lD��$Q|d!R�j�q��/ub.��:����#	��>���lw�o��Mi��xa,��-�ձ��s�
7E���Ƭ��	mH\^��*�S|�$��2�w�RJ���~H��<O|�a�x�?f�`�ͮ��f�a�Q�,���[�dDpA���:yz'�L#x�֖����֍�Z���#���V�/�i6^�v �;�n�Գ7l���N�L�����r2�eG�fl���'_?����� w��(n�Zv��_wS�-I�u��կ
Z���C���M�m�mGH�.)�p]���Ы���}:!G����lt�/�BG�~X`v�����i���u�9�^,?eoX*r�h�Q�K�=w6��Mgg�۩��|	�$�/�P��]Uш����Q�ތ6�-�	�0D��`�O�����vU��3�4>���̹m|�ڍic֐h$�?��*�@֓W1T8�	�����(��d�,�`iWΌ����AGT�Q؅���U[�lC�v��Iٸ��3�2��.�_]��pJ��^����Nt^'�,Rj�����*�>Lp^�0P�]��Sq��Mr�k��M��U��9��;nVI�}�~v�@���ǫ�Mb5��s���p�W$ن=s�х�F��OU�P��_*B����x�JhCE��M�(���ձ7v���5�$�/�?�^�r"���>���lO���zڔ~����������f���f�XX� 	�kE�,�-T���~EK9;������޾t+JTn<����ቂ6�*��`�_C~F9݇jD�tn�%T�a�����얋7��T8{*o�0��&��J�	=�/�N��a�}�KJ�
��x�ɨ"�7�0��tA�3���F���>�j���udR�P�ټ<
��P�QH��9��e��C�A�r.?`��D���O �Z5�J��K��S[��
˼]Z���p->-"	\��EA��</t��4�$��t�s��J��S�
}ѿ6x�ط|?������u�
��1&��B+�ҙ�	�`���ƕE��T�C\��*MF.f �G��%�JN���o��G����P�����^�C̜ڥHZi�Q:]�3���}M�7�zQU�ݲt ��dwv���	�	]��շ�|t��+-X�H�W�+��λ�I-�'ŏ1p�1�Z�� ��,#O��<��r������� y4hݎ%(iJ����`;p�&Nv&B9����n�^�כ֨{���/����N��+�]�d��|^��z���E�(LzZMżm�!�GB�x2�\M����O��'^4�U.ױj� �U�G�Iޛ�@V�o���.��d���@0m	/D�*��!�r'gK�F�6ooXW��-�[�U�ͻ��ʆ�c[RMb��ۗC���`T� }]'��@��#�����+�K�.�>�({Ѻ����~��)��,��X�V������̷���P���O ��B���Ur�����r�����)��ã8�m�^�bDF�Jz�Fn*)
���yv�Ij��	<]n�0�LWfhcTTP�ZB �G�'�eQ"&������K�l��o�Lx�^�Rk�"x�.n�K�\6���2��D�!	N�����bK8hm�+�o(��6k^H?�aR�}�I��e�D�4Q3zI��ʤj�0PDgƇ�c�d����/�hui�*r�I�.znܢ��)+?:�W<OjGz�`�{�P�Xr �)R��N}�Q��EҠr�I�|koi���p"b^��{�I��� ;%Q���Pg���ӑ,ly)����ޒ���{�%��i(����	e;Y��!i"�P
�����n��94d��|oD�(��W�����G�^p��|��H�����s~�?q�r��m٢�h/ <Tx<��XQ�eF�D��yM��?��ⓥ����瞜9R���>U�@�J�����4x�6�\���I-�'6�Ds�Z?%q�3����	�3-4�^����}����=�K
v��Z�bI�&��Y$^����P�9� nÁn�J6���L�q��`Ou��4"�2��i��_b��դ���R2�#K�y䰃ٰ�w���U���[��e���%7 r�<H�a��`s��f�����O�)��� э�Q�!��óٟ�8�iȗ�O��i��Mp��m��x>@�P%�����+�/��=�!8��R�X������\�H��H3�T���a���5o��h}�`J"~]N{0_��}U?u���DA[�f�`�������$��i��`��Ԗ�}��h�>���)~Iw�"{�W�k X���$�u�@�#|�-��~��=���2�^�����`O*��mN��8����x����%}�6�z���X�i����+&0Ӻ���x�/of6ei[�~�����P(^��[b`s��1�A �_�/^���35zL���"�^�kBo�Z���D�"�����yo�<1��h�9��5�u5�o�[���}��_�Z2F ��*�s6�$"T2����� 0:q��{�)��؄������X�y���ј^�����Cѣ�6�$�W�,�"����֛#���ꡦf������wQ�?��\��A@�˶f�+4
}ta����8���K8l����SW�� p
������͸��C�:�6�o�$h���^��Ǜ��6��Wxǖ򯝂O���F�?��F3�`��!��M��:���Y%�)Ů�.�����ބ_�ȶ���}��{������S�ZT�q��گ��C��4l^]�J17~b�=%F�xiF6@`y^Z�w���j���o��W��SA=V��;Rd�jZ�R�����NT.@�|�η�K���1v����G�]Q�RʘJ{���үBxM��2p�/����7St���7�J��(��+�A	ji�������Ti�T����"�n����@$<�L�d%/���p��Qf��TxE�?y��+��M3���Ƥ��Ar�扦����yn�)�8��V�Ku�k)*��-�|g���l�l7��iq�ϭ�.������x$^��:#�����s�	I��Śz�M's�׭4�)	��	�壘u�������TD��jyp�Ė��DȾa��I�ۜV0��_�y��!�/�&H�p�G�X"7�M��)�2űj.\�ع�LG�@�rw��6����("P�1�:Ź#(�N�h�q�X�~3�ɇ_�-�]Z�S|��&W2�Nރ3�!ްn�r��u�'B4E]�a ��[Z��GȔ��SMK5����f2T�;�&.��Ԣ�@�]�W�5!L��j�W�<�6�h�˼�Ã�1�ڨ@>���C��_׸�3�#=Z�[*H�����%t[łA�&:�p�)��=Z�e,�QݵwnNYz5����TA}ÂhcC�V� ���D;w��n�4�~�44i"P�`)�mWk�P�{_ ��%�u��{�8��H@�_�!���� z/ڻK%Q��ƻ�U%Ъt �F�Lң��i;�Z��ԾP]��ͻd��ZY�JU���;Uq �1��l�jUD �i꟝�����spw�:�YFh2����ir���� wB	_�,���R""��BG֌Цl��;�����)/:A�(�sfs�"��~��sy��*R0�'%���Va�᥉v�wNr5���@�@�b��*^Ω[u<�_�!���K����.�����̢~ƳA�7�KbӬh5�Y� �;ҙ1s���R��׽[T5x�GS�W?�ǝ��M��e�ܬ4:
VH�@�0�E���1<5���8L�b�w�O��b;n}A�l��㏧ʯ��E@��o��Pͯt�:��e��&5��s�>R�����������i����>�L=��j,�|��Z?l�?G�;���Fl��#��7-�/��0�o��
�ؿ
t�ߝ���m�2ӆc*w.�O=�ޥ�L9��"�h#�@����5�ԍ[��i#��ݕ1��j��/��Nٓr��: N-R$�UW���ƀrz��@ �M�ȳ"O����A�nE4} �,��<�ϛ�L�����D�M=��dg�f8a�ZA��G�h�>_����m�5F�1lv��i�V�n��$5�f�j 6�4H�A�/Ya�h!�9
�|�PKW���:���Ur^�_lfk�rB>!�����֞H���9x5p��e�2}���WN�n|�Z�q@D��Ғ�%]π���[A�D�9tH�����`?e[�5`R�
	��K5���u��V:��η:����U��"�VB[LW��)N����Uw�}��y��5+�X��.V��{Pr���S
hy�K*x
��G0D�<RB=� �t�!V&� 4|r�����>�Ozp�a�%h[lh��n�|��%:D�K=� ��~�B�Sps�;�b/�'v�S�CMw_2�H�cL�9]>)<�4Ї9����d�svg/!tHz�ZT2�@�u��\�M�9 �Ͱk���6�_�F4��&3��-�ff�U�v����4q�;��Z�w�F�h��h5t��ˢ�r1T����;J�Bp,�K�
%HՌՁ{��7�M�:Ď8H=�&i��6d�hD������',<v��@̕���lAK;�BړL��6�V�2Lc*fP�Ӗ���wm*]�B�J�E@{x�{#�����y�zC��O!��rd$.mz:���1a�J;)�Ձ��~Y0�����6�Lk't:���v�9�P�B�x��Oy<;���G��ҿ<�y�(i��:�C79��w��CL�<�$�"����cK`Dk����r
!V!�Ҕ2;��U$.m�K�^홦�9�s`�.�z��a��@�$��Ă��?�Qo8�p��]2�v�G�$��#)]\��Ql�@N��c/q.��x�?����v.d�i�M�+N�C3;���"��*g�e�Zv��z�!��*���B���Kp�h����v�+6٘�l?��}��.#&�ĠyQU9�	SX��I���+mD[�E��s�ڨ|i�e0�U�T	�a$�M�]�MG�1al�\�����V��v���Y���v�Qk�>�u��E=�v��W�?wgvZ'=�h��fH:1����4d����,�����=s��u������H�mqZj�oS@*��{���z�6ִ~ ���[K�]��������qn2��C�T-�Zsй��YW�J)�d��(%��mAt��S�%��5�'ٟKn^�c�:�?�5Y��k�s�W��E��t��\��<�b|�m�'�����4fb��E��9A���&Px+f�{&�$��e-�f���Ϩ��/<.&Lu�c�y�0Rr�E��tߥJ��'�x{�E�rMLS�i��Kh��x�x�O.p�aK�W�!���&�q��hπ����Zb�j�L�"0�����2vx/�ق�ǳ�m����Ɏ�6�X�@���'7�������YA]{�:xX�/z�oϣ-�mX����"�D��0'X�d��g�a��݃P��M�����`���$��:R��V�2A�&�xp�ɻ���A�T6r-���þ8 6b�@�w�Wm 1����Hʚm>+����4_���a����e(q��.�s/-�z��{qF�1�_��>7F(��&ޓ�ڹs��,�2|��E�t�
�u�,IQه�!�����IU:1$S�U�Ke¾��hB�� �̠S3[�Ы�hʟ9\��6��*�/�&���	x��Mx��;�?9��;X�K�CM�UumB
��/�����I>X&����g����M^Ws�4����<�������w{�]n?�0�7�8���DI)(�����s}���$���gk�F"j{@V�?�!,�A~t����"�O� �{���ڭ�-)8�^˜����
��.��_/��(N����՜	�AJ4Q�5�p�8(fa~�J K���4����"�9��3Cm2�[��8P����P�H��v_��0uc���`�R��:pd!Ҋ�X���'<�_���Ӄsq��m��W��}��嬷��r ����p�cb��<�]���9���qEޛ�f�#�,q�Cz��:��i7u$�����ն8�!P\`�xbƹBqO�`D@��;u�� ��W�	)��UT$���+O7��^�yx����Zs���׹ݷdg�d��ժ�ˣ����LM�,鳐�����8/)�\o>U_���S��`��k:kW���m�#M�Af����~l����UH2���;U
�������a�<�ߘ�ԾO����t25d�fBC��(��p��9�2U�D�I.�W��ND����\/�t�?OLk���aD̛���Z��=��j��R���Q�G�.��p�yt@�ЅI�Cq��^��i��h*,��HDC-��g�k��0�`�"=u�+�9x<�v�Z�2��R��vHXl��k.6;sT����b�w��6�2��!��P��^n�b�ۤ�R׻�<��$������PLY�W5(�9)?�ϧ���'�����i�{`�iZJ���Æ�Xvn����L�H6M[BA��} ���LJhJ'3��]֙S>U!��ٚ��1��lL~���������Z��H!�76mu�~Ӈ(�F���E��(M�tl���'w,��F�Th�[3����Zxx���a	�J��M�Ŭv��zjU��
�\����pާ�Yǆ|�D�\���)����x���+S�s�l�|�����y�h���:��L��xf�!��^��\��n���8牘�Is�@�v��c���v8E���,)�Y�1^=K�g�$அ+�NE�>� ���߮]ط���|b��G]w ���:���F�9SU���+�Q�*�%J��lK�OV���X��}��tIO���}��!f��Я[�g���ogb�j�{����+�R�0��kS�H���<ʮ��H�V?��qqa�6̄)*����ݱ����=t`�tO	�\��X�(8%�B2Oud����#�;�̆v%�9��/�@L��角�+֓qv^0<����ؼy����ja�Ne!�:�v���ziD8d��N���W�9�H�i���T�_���+p�[cZ�,����@�A�P6ɻT;�|s�4�%P�Ӯ6�a��t0N$f��M�0偼L�dg�ř��zJO�,�����0\[��,e@X��;[긚����MK���#�^�Q��ǣ�uc�'f��0|+�s7�Q�(�ԡ-���[`�4h1�^�C!��~���ޓF~��V#y�ޡ47�\��G��O?9�{���tM�^&nۃt��J �@�ܦK+�aZ8��`��˹<�'�o����5G�6��jH���s�89�7)Z���+�&Au�|��4�W��o�ݠ�W���)l�s�$�y����$Z�j?�P�Sj!±y��y��f�QJ��:HE�h��Q�T��x��;�A^1 U��h�H�I��mK��3����$�c������T�c=���;���J$,0/J�e�j��6��B%\� ���X������q)�}��΄W�U��&�Z����+�rϰ�w*��ؿߛGs�'�;!��G%Z�djk$6*A�2��a�N/ �ɺ'���4�B�;Ōe=�g��:���g.�AV�������~(J((@6�3?�`���p_vK�Zq�D�����+��Í��V�1�w29��wy$9ر��z�77��u/\#�v]@�S/Nf��
%�\�Ů��آ�jN��S�C����]3G�ʒj��֚�r��I}.��͘����%N�ӡ�D��͂id$�$@�YX�*�[3���](TS�X�ƖYw���)��kA