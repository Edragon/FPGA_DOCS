library verilog;
use verilog.vl_types.all;
entity and1 is
    port(
        y               : out    vl_logic;
        in1             : in     vl_logic
    );
end and1;
