��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n�,˪�nz)����Z86�mΔ>^�!:o4�\� ��n5�d_ ��s=��Z9&m�9��=���߳4k�a3!�DJlml�Z�8�d�0$�C���D��qU8^�϶�:P\�y�9�5���˂���H��A4%� �s�@F[�"BZ���=6��I�B����5*C��}�?+j1���s�y���HkeުA�%{���K�gJ��hV�o�r��'<99��ܭ����G��h5�˚�Vg��ƻ�^&���8�X���`�����p���5��#�(t��wuE�AB��%V�	
q�O޶T�d"�CG*�M���d�j�M7��6D��J���/<)W�j��(��#C_����|�$�5sA֦�����.��l\��&Z��}� 
����h橰�RsR�;����Q���F)��A禔y�!7M�}�x&�#r�hhʡ]X�8�E�k6`��?k������5���V�<����������C�V`�_�#�_;�,���y%F��e"�J֏�jߒQ���R���;t[��J�W��IÃ%�w�f����Њ�؂���B��x"k)�C6���i��9,�ЉeXA?����MM�,�39#�̄�/�^���6��ؠ��e�b��@j�#١����.������h��P/��"�K�p+R��M[؟��zI���X8t�7p������@I��X]C?����>����=	�U���������K�����k��Q����x���|��+�$��4�yގ��XA V,ʆ͗`ɓ2����Z���*��aم�hY���"�h�^4�����F����ot'Ր�](v$<�ʒH�W�F��jg��Rs5ٜ��S���)w�Jcb�$��=X�(��V�Rc�E#=�\m�*�ĩ��;wF5t�c�^��Ľ?C�;u���c�=7,:4霳��n\�2�Ȑ���*t�"'���6�����	,���2"Jm��邏5M zG�²O�B`�h �^r@l+��[���v,a�<|0�B3���Jp�����8g��J %�~�%˄,��Z��T�0��}�<5q����+�C��\3�aUH��Dn�d�m%I�?w%0m˿�O�ITmZ�i@�n���9��9uk�F$�@�UJ<aX�ήn�[U�b\Vd�i�z"v���WE*ǀ(�Y��h�n�OV��0Ww��C���b~�����x:���P�Xnu�ثn����o �I�>xԛ1�3��n{�HwJ I[~v��'Cv�Ղ�X�4�����R���X��/�O01�ՃK�Sg�,�FPh���e�A7*�F�SQޙ!��A��@���'�.E�b 6��O�|�yӔ��d�Bu�"�TH^N &�xD�VW���P��y��%v�э�3K��Vz�,�K�� IP��n��6L�u�
�ؔ]Ȑ�5kʋ����0C-'H�B�\��u���K���L�1��I�<��s9t8���@p��z]��F-P�*��3Nf���_�Z��� {|��qA���S�*�Ӑ�xN�x�-�_wY&5XlD�,(�x�.\�yB�v�K�M3��X.��ja�=�~:�51S�jg$韛���I��"�Q�H����o�k��e��)�XE�@��y�]&���ͽȖe5�J��:��*#�5 �mh��d!����!d�"�a�@}E�3Ov؜��o҆Wo���g2�tHLb��8c�L�ބ��#q@�U�N��, �@���z0*`�
�*5�q��e��M"ﮜ�M;�jy �E(l����0s�ͣ����ԫ]��4ʟX��,�@5���B�w (v��%�2mԾqW+?pV�F-�K���tÊ��X�0�Ha��&��kQ*^�������=t���t�H��vn·�E#;\+���j���b�S���:�V�D�aՃ	����\�nk� ��dH������'�zhH��'�ɿ������'���U@�-��|�}ꐪF4d��_�^�}�I8�G.�η�c��+����D�3q��_�#��#�Fc�!JX @f��ڍ	��1('ށ2�˓6����&%�x�k�����_R�'θE�zƘL���D;<����{���gX�}ۗ^O�N��gP�$+|�W�ڪ���6e��pe�FǘG۵V��͏���[+����l@	y��]�c��
�����ȑv��i?���4a��ߡ�x����P�$��ۮe�j���y�G㳭�돽�65�B<��R�e���^E��v���J�� �d�I��6�t8�$J����q�b�Z�:k�1~K�Nv��8��b���Hh�d*���A~��,�&��G�~;�����M������X���X ��9A2-��)@����w�v�Q��h#Ѯ$]X�jy�.+T��D鋣�tӥ�Ɓz��af��?��zF$����[$��8s#C�#J�A���L'Lx�:��y���k].��x�h�B�����!y���G2W�kf�}�sɦ�۱1�8���]���96C�j9ͥ��K*�=�o
�ʢT�k�C�"t}��T�%w�{C����Y���ZY���o���op��[���T�_�v�Ժ�_'D��Eu��x6�0O�"�ץ�Hm��rG߃�#.�;��ó�&���12/<��r(��T�QX1�g��J�Y�z�N1�aK>��"��<7��!�o4�T�)��p����5U@��f�%g"�����f���Tv	�(��W�	S����P�2��x�����R䀞羵r�.��<��s���	N�g����4�B?�h_���&��_�"��Û��<�aJ�'�Gdk�mw�4�ɘ X`��; rz�v%9N^u�x\�`=H��NR�J>�y#H�?�R�k������1�t�p�$�pڎ�S��2��~��p�G�������v��2�-+ze�&~��)��S �إ�K�+���^{})HF��|0N�Ҥ�r>�n@�J��E���y �FQ�-�R�
K'l� ���M�*gwƸ�g0#�DQ�z���9�-��	|,��ol�hwf�4nwI�=��mf;�0vJ[���b��B��:[)��#�p�l�����D�
�X���JjG�j�l�YGP�qgG�?�����j�0Tp���	���D�&�	�OcUvCq�i&�f����/k���\�dU�����Ӄ,�ۜ~�v�^�w�r��}�GR�+^,�����%$)������w*�.�0&�B�R2H��yj¬�x�����)��l9n�_ҝ|���b}��qEZ����7���c��e����T�q~�l���|�c! �����Y�qY���_�j�so6�t?˓��,H�Q�{w�]p;E �{���[vec�b6x����2���ѾM*Ձ��d�jŖ�m��F{i�;jK�:�&i}ۤ����k�fDo�����7"�y�	�5��r�p: ���
B/� �L�N��$���G��UCKhc��,���3��8K��b��E��+(����}ɊYZI�z��[�*�8�2a���l�p=yh & �b��d'֢���a2�p��E��%؋�W��S��~k��*��Z��-9���Q� :�����-c���_��!���䁳V,pyŰ��S	l8��c�٢d.�������!���.Q�z�����F]�%��װNӹ�����l������v?&�jJC�8�:%]��h~qQ=���!�>��C+�i�ڈ��(��w}[�p6<x�ۚ��~wkd(��r@��9+w��j�"y����B���[x����� �W�k�1�9��A�aa�fҨ9)�ж��`/l+y�JӜN��L��Z�;)He��R���y8pޅP�B`���\[����+ϧ���0!�d����{��a�)Y��v��7�(��D(�WE,:`ovD�{��Z�<4�$}$�{���������/��D���+d�"@�&e�w�5�.�k\�Y�����K�k,����}Vڛj�o�K4��\���C����Ap�����%�F�������P�X�����Z�y�<���z_h.KfUy�^�T����[u���#~�2�Z�Rj��[V`�i|�Y|Sbmd��d��b������ܙL� ��������3�;��OQÙ�oZ�=X��*�G6,�+3�9�O��l'T��K-��=�~p`=}���ߥ0����+Ա���G��עu�+h�T9�}D���$>U�mX�����;��=.q������� s`�-����]�&�:��[5C�Zo��y��S����a�Bu���h� >K`�D�٬��a�n8" d�7��Ѳm�D��eo��8[>�+)�.ۼ0��5ZާJ0dP��ު���]
����#��u�/LpW,�U'Q�׳X6Ս3�H��t�3m�:G������z��е��nU}~@>t������,�J~������Q8��Tz�!ėPu�(����%��u�b$��=��&��o��:T��O����!����BAz�wë�Ѝ�n�=�I;��s��/�����R:�wg3q�*Vq�ʭ�F���&x���규J�ܶB+�x<���y�����T�7)
�ܢ�'Oh�`�}~f�g
��J�)X���$�<�n�z&�M�n�Y;]�X��&������t,���%uj8�����f�g�a�9�d���?��;גA��!�}��<�N�?�HG��l&��<����+97W��a�3� $R�삗��I��'�tΚ:�������|%���8�U$���I��ڙ,,���nB��|*£T��n|�v�S��:*�)Y�F1ԄM�d��!qt�Ι���:$�}�}�������f[�����3u�=tȃ����<N�w�>�a6������.�b��l9���&c>�'=Ͼ'*F)�a׬͛�^�\���exq��RW�	u� �l��)��ی�.�-u��j��N:}qgS��#N�'��壘.���]�%��6MM��Qq�tzh����2�|m@G�;)�̈��}�rzS�R�^�Y��=_��ͦ�7�k-`��9�6���i�Έż��۷\Mq%*�v!l$k�ً%җ��$�?J	$s�ؒ1���+O�%Ē����Y�#p}�D4� �;eH�����#��l7\K?��)��X&�1i��1'bԃ���d0e3�p�"�'>eX��FQ���N����^rm���Њ��Jl��F	��C��1%�|�q�p�Xk�\�a��l���t�N����\a�ۼ:�_ b������,�p�o[[��uvs+��n�Z���
��#o���L!(��
PחT�c;���ɜ���<�i*қ0r�Ϫ�E���n�)}%�����-�e��D�4�3����K�d�-s.�4 ���|�-�w3g�~��B���f��rНK�骆&��K���Ғһ��O�e�Lg�� �.pj!Uk!�a�вำ!�s7x
�3ry�����,��(nAb�\(`��Z$��5�[�rrźl<�%˜�M5���-�U4�İ7��Q��d�%��Q;WS+:�P���w54�Xw�PO��.P�0���{��|ڇ�]�JzX��!�,�jk+��pF�9���� %���Djz��kc��L��x���]�`���X�7��!�}7��|�Z<���Q]8��&P�(�%W�;^����Uˊ1�W�$�0)Y� 