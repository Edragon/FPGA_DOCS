��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=/�b�2uM[tڄrq��-�{N�s�p��U�n������L������sQ�{_60+y��g��k��©��Z������<b�)��0[8�:�r�Ԓ])�Vl�+R�}�cD�=��wR2�ũ-Ij�X��	龼��u�������B? ҕ�01�6�����U;���B� �gt/`��V�:w)�B���Q�X{�ޭ����bd9c�o�aɒ��S��x��<�5���C�1ݸvK���
���v0�$�����nv\�T�8�.W����)��Y�|_��L�{ߓ�+[��5��K��/(��JuF��#.Kr�4V���7(�Cn�	��� C�����2�4�Hռ���̧�4V�x��*p�@�WL5��[�K�3�hW��F4�Ѿ׮v��ii�d��n,Z5e��e�/�g1/��N�8òP�׃���E�~=�������G��s�ӱ��|_0�\cS��*`�0p� �5����S��_��>��)ɊĹ�����ᝈG�>�ƴF���Y�w�'�a�$@�rY[a�+�
Ǹgt��.�)z�+�R�{|�����>�@��֩��J�)��P���YR5H���W�]k��/�q�Wp�w�p��� #ef��>:�J-DKf�=C����-�.&���;��\�����56t�����0���R���x$A����^㫲�Ū����4X"BL9�6yT�ʏ�3�?B��&!�I�a[X��w� �����(��5���[I�[C� �����m�
v���<�/>�}�� �����m��%ɴ��-�FZG����Z�6t�_b����b����=��r�Su�{(ؽeLC�ˉ�mm�k�L�kho�N��Y�6���8�g�ɫb-��B`�Vcޑ!�o���@�����i�-���#aw�Gݩ�W�o`'eP:˷�6U��!�����kw ����?��EʔI�m���v��F��J�v���6���Te��<b4�Wf�:E�P���~��NK�{�_ ��P0y49���K�y`6n'��_J�#M|�z!�� <s�������R�謹�� 5gԲdO���N�pf�T,�pjƧ�,�j&س���-���S&2� ��@C����H�PW��B��̫�����y�����!+������mY#�x���zgl'dP	Z�f�bθ A���ڪ��坐���&N�j-؈�1������9�<g[�=��~�3��r���R@=Kc"j�ܤRA�<���U����P�,�4�������k�� *��N��^@��3��Z�M�q,�J!�M��@�J�μ�HoR)N���	,7�����"ԕ�mU��E���#�.��K�"-.�W(����8o5*td��4��n8�cp=�C見]:��w�&�9b�[��7h�E�1�����^�w`1�f�B�Ũ9.��1n�z�pߊ&�)C`l�%���rD��N.d�@�:�_0te�k4��^�Dǵ�吔���>/�6�t7D�ٷ�_�Xf�r�W�mԨ(=�ɍ�&�5I�D�O�{k���&�"k�q��%����R�K���O��L�th�6;Ǘ�<�i��0�(m�C�o�J�n����|z��1�A���r��w
�*|T�v�р�'��'>7���e_Էd��:H<�GJ�i��i��`�]��M��J�h�p��C���"���9J���H�]";��y=�>��_��UWJ�����Kߓ�Ÿi���d\���(�)��BZ�!�Ț��᾽Læ5l��ߙW�9[�+�A��1�$A���dn!�H7&k~�J|�Z����:0p�t��\2�|a㎧�f�o��s�g��I��N1� fg�2|�Nx��C��U3�,k9�u�$sֱo4�6�7�Xε�d��;���7+/�輚T��aU��9�j\���J+1�#9�o���� #�i)���}o��γ"x�>�x�q��W
0c �\ő/���,K%�8m�ph�K8_2�����NP�*UE㠈H�+����dw��Nf{JH!	z���/�I�
��Is=3��}�$2J���^�E�����@"�eA�u�w> �~����K8�dN�٠�'����D�#�����m��s[�ۉ��~y�?�4�W�,Q!{�[�g�sx�\�=�ڊͰ\����n��	�^����r���K�R�^{�2-ydwǬ���zA�1w���x9<��b ��	Ի8����#���"�Q��+�=s���3���"s4�>��J����+x{��7�y@��},�s�B�XA�e_��>�H�;3A�W4%��G�\���&-hD�hGi��ĝ�b%hrᳬ���&�H�h���v�����Z�#��,v�2�2:݌%�wL�lthZg�6.���ϭ�32�7�����\U��2ÁAk��H���I�DSP@&�<9@uCc�#aDH�KA���h����Em7���G�D����R�^x�>�X��6����ä\�+*eP"�Q:��KЪUGN�UZ����Cm�L�W UP�} ��g�!���O�oQ١/�zد�8� �r�� �zª�d,����Z]�ډ�(J��.O����s���)��Qh��Y9pk�^�i�C_k-v�zH��R>�w~E)�u��B�H��a���%T�\�1i���	f�Щ5k�l�<V�k��qI��P�2CFy�˺.�Evt��J7�F�5efb�J�h;�����:)�h-L��>�}���:-��M���^_3�f�u�"xQ�{��U8��*��E��1^_��9q�œ<A����ҁ��ؾ:@3t+������ʿ���ihYh������ˢ�2��0H0�"��Y�/�#Q�eTHM��|ZSv�,a�}�!k����̪c��>���YJqb��f���9.S�}C2����^;���5^Ш�fhB�S�9�In�F��i�<es)���La���5r�%�g�JR��{I�im�uP,�D�Y�;Cb}ͺѾ���DD�OQXC1g�0>��Σ�:o3	w�UZ�IΌAS�w+�}����n:_h�C�y梺8��Y��~*Qbl@�)�7�L�
�s00*)d��ކ��p��Cm����ox�q�d���^#��x�������? �_�a�r�S[����l0r���/�h@�B��a��4�[O���3{L�=>չ��+l��յ�d��:x������37�u1��5��yX���> �Tb��E��dt1؈/j�����֖��IdA/Y{�.7���vg�ʥ��g��<,UI{��w���o�Q�m"�_$�9��A��u�BYg��j���Y)9%^�,�I�nt�5�1��M�m�BI)�6��~
i|de
-���� Ut�~g젨�(y�1$�ⱨ~k���&�3��.�RS	�L�8�d��A�7�N����Z�r����z�E�����
}o���w-��X�0�	�sF���A �Z(>Æ��V�_� td�t0�bqd��҅Yާ�EV�ue�0�]I������g�?zD�Y1����U�{lQmVy���/�k&⸚U
4�7@:&��(�ʔ��)���沮� KN4O�c愁¤|��"]+g�.�)�_]��v��F�ox�Gŕ���|�-z�^�|L�2Q�-*t�nuض-_>nx���ef��Gk���L'%������,�f�$�|ە,d�iL�o<w�cYKt�^)a�_X.�i���J�0i�n�BB���=�`2�Aǣ^�cJ|��+�kCz��%�Bqv�9����U��Q�$��lr8���^��I��v�qέ6(�Y����a��F��T�H���q�N�e��I��S�o�;�g ׽Q.�܆c��%+LC�-�qWOn���V�!��X�-�,'��uT�@��gץ��b}�#�*����O�T��gOT&*�� ��\ul���rG�!��!�(����_M��B��ǁ��<I��V �)�e��f�N݅6���pZ�C�k���M=��u��`4eA�h�-�@p���$9G=�c�,�A�=쎒l�6��A�$�L1ł�Fg� d�΂���+�Ԧ�M6��tb�d��|�P��2�������&]��/F.˘_h$�Q���nFbQ�n��
d��p�"r��J�B��К�j,Կӕ�!��D]�RlTF��M�'żve���m"� ���i*��
����Ҡk����w���>��${ �5.l� J���F𴬏'r�[W��F��������i�Ǖ�
\��o�za��+�/���s��C��݋B4 �R�T��{⻿�s*��<��62G"c��^�fr8%�y�K�r���j�_�'��=��-<�c>$[��j���� �u�e�;����z4=,��@�Ld.��K��4�:�WI:K+����KJ�m|�J����o6����I��KP�-r�d�k��i���-ta$����9��1�q3ثO����K��O�[��ݲ��?�(i�;>���݀��8����7/��%�G�-u����@P���)�_�u���Ѱ���ni!�s6�9������
8x�����3kMH�������,b<��(@���ϋ�Ptͫ]b�f(�L1�kX�kE�bM�	��1���)㋋%����*/*�U�/\��E��cD=J�SaH����T�C�kh\Ѧ����3��ךd�J���H�rЮ��*�R�؂�q7+j�@;��cG��;�[�څM�Q����H7��F�0�&5��ʧ��&q�b���՚��Ĝ��!���s>�0-<�x��GJ��vH�D$��-Yu!w���I�X���"[<���*G���`�����!��[.ƌ�?���i��ϐ*{�sɶh�z�,|����ɊB�J)�ú�+���G�c8������p35������e9Y�Vⴏ���$%%%N�ۮ�)���!/�(�s����H6\��'��ͼ�~����m����y+e?�\+��;��&�8g����14���&w��o^���ת1�M�+f=o��g�a�m�Ma�P)1�T����/�\�r-�1ܘ����Yy��\�����g����V~��:�o����5U�9�ܹ!�No6�7pTX�Zڭ��Bm�۶��O�M�������C��n�����)��+'}R��#.m�q�������r`�:Zz�	�A�b���\��,��k+a_
���/:fx�]���5&�I�O�x&����k#K�1�m�.^�c>q�^�(ƣ%��5Vʻ�^���Hu���H�e;��>����![u�$f�̅ɦ��a�|_���D����x���u�3�,����"��Z��(�w#EϷ'<��N"h���B����\S#Uhz�+�sfV�$�n�',�� J���GHc���*��F�.��<�	���r�!�e;O;��Y	L�����6�H�3�C2�e��ߙ�������<I��fS]�!ףr=��%+Y�J�hK�BZ������N�ӄ�w�Y�fCW�S]�6Y;Xpа~�	��O�b�N���y����tT���EKSQ-z�u-2[��,�>/������#E\Q _�3�n��0`�����8+L��[����7#��}`���$�:7[��2wO�T8�(��_ݨ�mj��n �d�E�W	�
+_����__�&o���X�
��s��T�g�5������^P�)[�`܅�s2�5x�w��ؾ���4�il����T��X�lx�s1�Q��2�8:���*�5��1�=�7=�zޚ	��'"�� '��jj����֍��h�Դ4�xI�\�Z�Zt!U�Z�m̖�;�a�FcL��aт��;P��m�;��3�0�$x��!�R9��	I��~]3/`��;��!lb~�
���ڿ!�Qs��v��Q�k}F�J|f��yЗ���_"٣H�v��ĔN��S@n��1�^�}�)�aO5N]��s�����щi�%8���"9�饞8H7f!�6X,⪊A��8����2��P�3~��Xڋ���;r<�!,w�N��7[�&�R�^���lh9b����S�}�%g!-gm�(����P��+�3� )�.�{��J��1f�踝�����>p1d��BTѨՐ&��#i����~��ӏ����Ƒa�i��q'�� ����
�9�`�:���j2�I������ߕ�"݊3h7YKʆ�@0K|�r5�O� Ы苛��9���&�
�S�`g@a�݂`��m�R��{�m�1Cx�R�5�2�=���1�+�[���(�cM�f�8�s�'5�+�y�,S���a��6ų��:)HS`���$4���3���}Gɸў���4R����W�^A*��U�-i��������5����p&���x(�۲)�Qا��ە��%?�k��3�Q��Wj��f��\��-ױ��@Ų�$�
n�LЮ Q��*��b-��;�f��U=�����Tс#bɍ��Hp�e�*Zr�����7�7���E�2% D!�(ب�3V�*hg����L@��ܔ��(�K��M{����2��mx
9�XR�w��)�k���כ�%�	��2������ѷ��\h�Z+�n."wX2�]��vK�#�CS/�$�L�󊆻~K�/��=�o�<z3Z"C�Ӄ,ȼ�Jrl������>�m<������Z�y��=�Y�JO�v�<����۲S��-�����+9�����m��<�ǚxe�JW�a$���|�|첒$���m!���p�d_W\D�+�(�9d�+�k�q�f7�:�vmŷ}:�� ��2��섟�7�zD��v�7��C�+Nj��*�59�A�����ᵟ I�z���%`�l�����0�^��M��cK��/@Z��l(��L���E=/��.vW�Jw�[��IjIW�iw;�n�UZ��a���\�ζ���d��@߼��)Ë�9FF��[��9�eP�H������h�F�·&�4���7��+0��x�M܌BX�?G6�ܢ���_�!h�V�1v0BSqL1i�xI��ї�D�N��Յ���T����W~�b(�Ntիi[>��������급�7�g*S��3�5���#�����ٛOϮڝ�" ��e���0�iL�܇���>4D`�Qg�Z"����|{�SP����?�	�g�ԣ ���J$_�Q�1�j�ol�y�cwޡ�?��=A�R,��h�hBiKj�]~|��Q����aD��51� v}�0gaorrsߜl_�]����,�=�v58�_�+��ߌ�MK�Q�z�1
Y�pG�^X&8�����ɰA!�	�y���?k���
�A^3A��X{���)g\��U5͝N��"��ЭXa��d�4��;�7�XRb�;���w8"(�q	c��6]��,�Y���g�ƚk�|I�p
�b2�����!�K��`�ʠ��;��dE����K��)�����J7��%8
�O9X�D�D�T5��^&l��<��9�8=�����T�H�v"��G��)�P��N۷ �U^N�ƭ��K1�"�� �z*;�Z�������޹iFf�5����,��:Qɋ���J!r��������Yu� !��=yǞ�T����3��ԁ\��Er�u��d倌p���)�a�D��'�A6���.߬/�Q�֙�p[�\ɝ�"f��� vUq-��A�|tg�K����Fa�7�������;����K�ɖƿ���0���#�THk��]��Ҍ�j{�4��7���!�E�������;�/�ő�	p��R�^](�
|m��)�&�%0�i�r]�8�_>�Gn��uF�ri �xR��ٮ"�N]�%E�0K��(5�׬�@,��J�~��O�	�M�e�o˖f-�]�Q���tB��ɝ<��_uFo�P�|qjF�}N'|�u� Av��R� �f��x�.���!⋆Y咏"���e�=}����76Z|w.��J���k`U����e�J�l���@&4��3���U�%��|���N�>�S>�f~x�B��u��:Tay$fA�����f0���W������*�2L�-m��n�^�%��IO
X�h���E���<�M��RF��4"�gˢ̭�i�V�qy(*c�yNb�{s�E�<~l�E���%�%�.'�fT��sT��j[&�����!a],e���r`�(��b�L�������R�4����;'?Vi�\�BE�k���N��9�)�ʹc�8��Ȁ�I��]��z�O�F�;c��)S
����Ia=OK�'�t,�Dзf�Q��H�Gζ��fC�]������x��a�*���B��\{<�ZZImc��X�W��?��Y�� ��Q��Y8=��v���_=�g���Z�>4�C��=��`z�yP�G���&�nE��=��S�y��	�m
C�2M���U_H��:�3ך�+��ԣR� ��U0������e�׃^�
�O'��YE8��cD���<��$N)|�J�0\�N����fZT*���3�T���7���u����6z4FuU��B"��7]��6�mѣ�� @d���p
N��]���r��h���x�l��ݖ�|S	ȹ	��-��V�Oc�cp����"hZُ����˨'��5�r�t=�<��$2gׄw�.�A�!N�H�Hە����Ԟ�[Jz���
�O�	gk=���m8�z�O���Q�TR�38�:l�b���h3M-�|���;��H��t���!�3�p4!��"��[�C K/�C��FK����L��%3]�䱵�>S�Hr%
��$F��-̟�	7�6v�7����c�����n�;�^1�1$j2���)���W���#�mb���h���`��{f��� ����D�
�U��4f�DP�ph�r���'ˬ)$�	î0��ՆuCݑ���:��l�U4Zh�|tH�����!н��i�n��K���93��jEJW�&srO;����`�y��� ��2ǂ`� �S7���:����<Y0Ω�wW� ���?�q�"�����c��D��d��"��	�Ľ�@u�q�F�msHj+�!*����㺺��NJn*�NrQ:U�V�QX"XJ�Fp�Ա�\Ñ��Y2� ص8a�Qr;�#m9�~/�]�ӱ�߱��[���Pم��E��ə�ɩ��#6P�(U�; Uz��ep�v���u���?�;K)�(t��G��pq��3G��2���WƆ��2��ڥ����a� �l� ҷ��e�%�;O�>/ځ�?�������nK�-/���;�&��no{���/#7n��b�X4[G�]�	�Ю��gk����M��!Ɍ��sai�L�-�
��	A�$� @��qLζ�M�������	6������6q?RW)����96kw��A��^^Fl��GD�]%r�@��UO�ĊT�����q�Y� ����<��I�A��Lm���e�q�q�h���7�5�VY�3�v*�$�m�؊�w�����ǖ�խbc���E���$�6Jb�b��?�f��X

	�1������K�T���	�y������L��gt���/T��2�Ic���-όAE�TW$��N�D�i'p��M̓.ʳ���0d��ߊz-ĐVtĵ���$Ò/�	wd���&�@D�"�;��]t(b*���AH�����|�Ԇ�g��vwO���D:���[,�H)�e~�C�J�>����v�]��b���mq����ut��{oG����� A�����:D4�D<`Q(�~�X��%2IY�p�i��a�+�����f�p_zd5E�� <��C�̣ݟ.d�VG�A0L��d(�^��$���(k]�n��b"���8�7\qB���g��4SH����}����a'����>�|��F���k�{���N�O6Du1�N)��s���Å�q�|�`�ek�-�T�H˵Z�!]KO�X���y�ySJzH9���u/�t����P\ʡ&W��6[�Q,.8�����XP��|Dh7�
-�o��.��=[Ne��*�*�=xi�d]H<��n\?U	�a@�H���P����i
#O̧�$�bd��d�]\�a⑪W�;����
޹���D����D���2h���3>��,~Udm�p�2�嬚�s��5�U6A�Q����eJa*��U���؃����#�k�͚��~V���5��*��8@&T�.rΚ�q��wk���,������i���Í�y;��`s�.br�u�}jbM��GD�'(s���}h��A'Gx��:���-�}2o:����&�����O̓��0�FP;���z�ڦ�bN(~��Y_;��`�Z�lO4]�r! ���٠�P3��Y:�ae@i�<����l������tI��Dq�^ʝ4]]Ҍ����oI�>R�_����ˮ:I�u9}tHm��5\�ɀ���t�""������Rͳ�p�\�J�`!��tI��X��!/�`�����$���["��d��+ܪ�� O�I<���g\�<c4km�5�F}�������ނ���i�6~�Dq��w\軧2v��Ih�u����p�K��|k{ݼ������V���A��������)4��<皛��C7n��/]�����D;(�\Zc`U?{���賈����u'徂�6sQ�G�{qyw��Y�-���\�8��S������^~����f4�ؘT����w�T�ZYh��B����>|�X�2�\�^y�iތ��-�B����d����v��X��D�Ҟլ
�5rCO�g�M��:V* �H�"�]J<����_x��}dxj��n��1��c�^ɺ�;�Ti����6x:@H����t�N^<���h�%��ϵ��azԀ������v��|�x�u)涃G��{\�ο_�	�g�FRrg(��5��|�[Fd��Y}~nk�A��sHʴ|�?�k��r�q�9_�ȶar�lT�S�Ay�aJ˔��<Y�c�b�_���#x~T�?c�մ�~�H���5��;Ҙe���E[�<KJ����[ ��ձ��RFsl��'��V}'��S�k���wa >U*�uΛ4��μy�(�{J(��O�����x�M��A~�B���bc��M[R��(ڤ��\f>�B�O=��ж^�75F&V��$'h�7�U�T�'�5K��'Ym������t�Ynh��7�y����bau����<�=��P�З��Ӝ8{p֍`6
�9S��/�p���5�	���1�r$p542vul�K)����w��Z��V!�ڽ�Ojga5۝�f.V7�����c?+�Եu��m����Q<����+��Q�_��N�	��ˮiݭ���̸~e�s`Pcf��uz�)"��n�P������V��>?/� ��])	u�G`�^/�H��a����u/9������V���a�-I�c@�U�ᚺs����P]nRo���إ��_j�ҳu	vV���o;�;diӏE(���$�<�� �U 9��e���i[ȡ}�"������p��
����?��i���ze�5K�M��r����O2"{�12z�z�ݬ�-ж�O����G�7Db�a�!�y��;�������;��h�`$����ؒ�d`�t�6��eV��%K/�q��#X�ׁ.NX	��y
��,;��ܺ�"]q'�Z>s�!x����'P�~�Z+�\/���Ka�LF�j��l⍈�	Ǧ�>O��Y�c�.�q��U�iQ1V�L�u]c�'O+��<x�w���&V+��m7���u�f�<h�wFO��"�G�rC�O��o��h��T%}��Yf3S#�)��:9���Ӡ����1[-�5��"�#4{���FB\ݛR�ms��9~�ʳrk�#&G͜��f�w�������ܜN��Ȋ��[e?� l���f����+�� ��믵S�;Ttb���Ŷ�,~T�2��|�܈xz�H�j��ڙ�#ύ� �W��F���iW�]*�h����$�S���c �jФ:M��,}�cq��E~f��Mض�����ݟ�	���P1��
rZ+�,I�}���S������}�XU�Go�5��(<���DxQ'1��d�V�Y��J
pr�$�T��:����;. a4k�1Ls]�ȓJA��,���[�+�Ye�%�δ���ό@���h��Z�����@��vjӆ0E����r%��pu��c���~pZ�l褚"`�~����;Os��8P��@�l�M4R�3�� u�e#v�ðoƸ��";T��Ѵ ꐈ�<���l�����X��v����ea����>-�n�1`�%�`n5e�� ���q��T�r���cW?�Ϭ	6�4�.�9[�+�u^���4@�-i������c����Ԁ1pzVr�ድ�en�N�-W��m2��7	�}^���Us����9x?*�;�1��pn����]���6p��?� ���[��[�w#�S���ծ֤�#*Z�)bulŎ�4I��ch�LY]kQ�H�^��%&���ߗ$���pn���(��6���-9�&�}3:R���d�\�	3W������KġQѻ~���y����g���3.�Y�ﱐjgp&��^����L�)˷���c��!�5[į�dXX��8r jڱ����!�GH}��EOV	��M씱;����ۭ�͞��D��G4�5�[9�6U'��/�
�~ì�˾�(���z=��#1U�r�@�ICջI��ȅ�@�TE� ��KCO
i>��8m
�(g�:������������K���K��:B c�_��NC����;�,D�������Q�h�X�m�=�x�W���4C��!`Lt��O)����E����Y�%B�f7�F\�9\{����2���:֓K��9Kg4�5q�TD��{�r,i���j��� ��]��1qF^����~�2�43c`���^����^�!L΀Z`�C���c�dC7B�|Сκh�.�RE��<;vh~���L����R�;g=�� +fŹgY���QP�dXr��b#/��c��Vz���#�%!ڢ���� �C��v��s=�`g�a�X��4�����F�����2�K�殌��J��/�\ �{|���X�P��3p��%��Y�o��_<�TC�Ft��.�;|�F�ѷ��*ϟ�o�Ѓ��h�e���4��г+n�3�w�=�)�}�����Ǽf�
a�Qn�XV���w�Avܯ4j��)D�>��[��z�����C�G�������Q�vK$�%�$ms�s����l68�͍LGa�[Y���1%#q�eq}�C��Y�m�ԑr���L# `���`#�X/�j�Q�Tw�~�?�:�7�͞:K���2Թ���\W@:т��c\���N��!���'�����c]��2��=�����\��OQ����RGp'R��c8���xO
-rڔ���O�-,S���B�#��R�޺3�m%ك)���<��&0t�LA��|��2��>����9�ug<G.
8��_$���_���
	q�'.���@�M��_\���
�ɐA�m�q����@a��4�M�h���������d�_y	�O�C��TY[����Z���@��sHR�c��4Κ�n���-�K����� �N^�1�r�t��/l�C|Q�ܸ/=�����h�,<u�jbj~��*D�,�6�R�~�,���e��q�N�fmЬ��A Q�Ւ�~-�f�l�Їͪ�ntZ K�t B��F���"[�d���T� ~�'M�a)j�¹��˖����@ij@����Re&�\`7�g&��6#�Y�����t(@"&-1��3��S���2�(������8�`���QLX���ٖK�ј|&��'�Pr���~&�͸�� �_�}G��%�w�7m$J"���z2byq�̻2��L�5�R�����
7����7b9�1�<?A`L��H导?�Z�|��#>��ۗ��.~w5��EZf��+1�u��1Ϝ�I�6�9Da�.��k;i�vx��-n�.)��Һ~��uOX���,wn���Lz�����N��W	&)��R �?a��D)K�
-��k>z"~0'�����S��F�=myƁ�?ogBS�0����&l�{����;�:�
,0�/m�?��YЁ�&�wP>��5�K���c1$ɵg��2�;�<(k��Nl�QAVf|�u��L4�G����>�<K^0��~���،[FZ��_���2���-f"�w��)�n$��C��PGX�A>�S�I&|��1HXeM�5r?�a"Z�6 ��Jgu�"�R� �|��f�4�Cb��kJygf�NzU�u\]ռ���5�&i�N2�̪�Ƽ��؅}c�Y�<�'��yF;��R�p���8x����уG$؝T���.n� ��&���+U��9N�N�rmo������'�@�f�3�DG��E��弉����3�||f2���������ͼH����JU�2�z�T�.lR�n؀�Ƥ�^���篿,��@��V�W	�/��r����{v���ǅ�/<�^�yv�.$�V��a{��Jn�A�Î��.����e�vVI�z��bw��֡(�y'��FVŤ��.����;S2ˣ�5���3�����)��Rff��$��<[Ƃ@骺_�c����]#��0} Cj ��k��쁟3#�>�������Lt�ycF흍�s[�y�6�Xǖm,�2��{�9ύ��� �$�f�ګ!�s]4V_���B)2�r��c�<��yZEX;�y����u>�̧�������h)�d�z�#����}��a :0+U���b�U�D���<A 0��r��	��P7'�^��E���W�#�Er���Dm%�Y�Q�7t�с��a���#5nZq����u9�6�@�s���>'����b�T�eD��h��`�2��N'O�MN!~���$W�������T���M�>�PD7�2�v#��!��>a�%8������*<8�?402$�ѷ��3��b%T���wR`h��d��=���w� ����Dal��P����~����"�L�g���W+"^^OT�~@n��;��&*RE��HJ�W����d7Nw�J)4-`���SS�x�W^��\�&�� +x��( bvGh�~u.ŖX�	e>C2�����0�fwPK���z���m4�G�x�F�ti�.̭E$[=��o��ѹOl�����ɱ9���v
��e�/sF ��}����ה%�T쟉g��'[v��w��M6&؞��?|\��~���5�*���<JO[��t�M�K9�c߅�FE��m}�2�Iff���L<�m�z��"P0ok��I �o���|h�xEw��K
�DqIsyK
�#vIG"�DD����LR�5���)�/���,���LY��DL�{�D��Wtup5�6���%��>��91�:1��h�Z�rF�7Ǉ�i���@t�K!�w�Zi��UO�sPax��	 ǻ+�!�:y�Ѹ���f�<�g�|IvC5�=]=�W�Nqt%A�r��4#4�E�l�Uo�����������#g$߹�s�5���r?^�h T�Ή@��< �+Tf|��Fy�2�[)�uZ�������u�y�a�����;�W�A�k"tkᙊ�TM�IF-w��ȔM��{e��=�8Pg(,����&����9������CQ]ޢ�">���E�u01VW8�c"����
������hf�n��.��,pf��&�A_�D.���_���o��
�{��V�x2��Cv��#%��VYZ�:��1��Y���)�T/���@������&/I�۝��c�� ��#����T�==�g�w��� c��b�z�Ye�E٤�1��UIX~������(��K�3zևoo~���d�=;������+��)���K?xt����|)�+��'������n�)UY5+;�cr�t|p�����O��$'J����PbȂ<�#�w��sB�����&����3)X��A�/���u��q��aB���<O�N�[�Z�8|S�~Ȥ�N[���`.i���C��u3�G�n�a��ާ&ו��z��O4T�4-��q`�5�oV��5YUnA�O��N�#��"i�!j}�@����]���kh�L�sF(�p��B��`�UU8B+�W}�$P�t_��k�-��<��B�4a[w��n�XbUK$ĭ�!G�y�L⿕Y�RԈ�<ڥ?h�mk������\H�����*Y=���u>H��H�*��g~)'I�y�<����"l��[��%���W*����` 'V�����)0É���X>�����]i)Ǝ��̷����Eg��[[���i&oֱ�j�-'"iJ��ъC�/-C�-RZn}meS�?��\s}0Z�T�������/��Tz9���ɻ��-E����C�/�q;�3vM��Z�5O���w3ɘ����d����Q:̺�?�,��X�<r-?=�-��],���5��1q+���Q��u�⍐A���D1��JK<���:�ˀA�u<��Y.)��Sxm��$&��p�C#��x2�@YƗ��`�>qe৾�/d�!���G7Z��x�������	N5)�V�n�RE����8?���A�̽B�i4��/I�۔���7�V3kS:8Y��n5�����GE��&EsK²bE�0ȴ��]�'7*�#�T{��V��I:{_�.,s��|3���nX>�
 �k���Q<Lr��O���eI���y,P���=�m��\8��xd��������y�����r2/��a�C26,�;1���Z=������;i̐�pU����ܠe.<�2��!e��ވF�Q�e�z�!#�Q>�)�Mtw=�-�P�G��Uu\c���X #���9PA'���Y)��:���I�����O�Ԅ�C��0(�HL-�L:�� �����`�¾�p�h����xn�3`�^�7��]7�2�ڽ� �=}s�e{(��7�IM��e��X=6Q�k��~l�ˬ��v�
�R�Kɬ��R�����3���JY]D��bE��E���U�[�r���H�Ҟ����4���H�B!(Y��j���:4�^I��d+w��h>���wf4d�a�f8SSZ�=�f>�R��&��I>�D)��H��P�p��eˤj"~@��-�m�;�[ d!����I�*����w�ͨ�5�4�l�ͤ����d�7i���t��3��:ٟ��e�8����ZC�(��&���r3�į�q�j~�W_i3��d�RN8���k�>HDy������������^����'�vJ�3O�I��n��!:�7q'�C���9����et��ur��������W�o7�q�;}@��3�i�}7�Յ�ξ��� BR�6��?LP�ˈ��iO$`H�����m����:����㶳O]`]��Dh�Y�ֳ�$v�L�$���x���
���<��j:9$�r5`t:"���VML�G%��!A	����"}WM2Ē�R���VnY!Ku�
+h���Y�RȎRiZ�QT�37��/2��-P�Qm��q��qb}�(|h�9�2�;�Gm�
��w[Û*�4��9R���O+[����p%��m\�F���U�(p����5r׋.~2L��57��?�`炔� ��V)l)�
�U�B�'QW��u��I����G���ka�E.��y�ݾ�ț�7�6 ��R���p7��^���u�z�Z�A|�r��o�� a
F\����B-E��7��5A�s��Ls���_ �ۂ����Q�q������'�)3������3��n4��R+�[ӉIx/����n��bf��"�7�׊j	��� ���<7��_Ԭ|~����`V�t��$��f��Pk���h���ƭ�O9�2g��B7�/_����PN� i�����s�Qy?L��w0 Ha���s���q��7;V�*�]a�����}��H%�G���&
��"V5�Ù�KQQp�Sg�3x�Jn��|���hF^�o�AӶ��ܺ�L���S��8�Ǘ�#
Q�ct��lhs�ܚ��0I�~�K�/�c*c@��7c�k�p�I\�>,�~��}Ȑ� .X����=��ƓbF)���)Br��pL+*�VP-��;O�@�)�G���@�9zmS�o�뻖��m�kc�;	��6���㪟�|�d����Ơ�Ĥ�J�*A�{�#+��m��1��_��5MK�����S�8���h*<��� W�;&~��xrZ/��Z�g��r�{�	�w������R"���us���A���u���]�5������݃���)V^�`���Ő_(�wA2ץ y=lEӮuz�褢�TC&3�
kX�d�����fX� �ɽ,7o2�}�WEwq�8.������	5T������@��3%(H�\��J�*���^!Y�'��W�=��R����b�k����8�\��a�\1]��m]؉�rd�(��/�`�2���r�k�����y(=��sadK�����[� C�w[P�k�lՙZ�o�&��{�I���]�B���*�|N ?�`t"fE�v[g#`v9f�`q�g�ϭ�_�W���ɣ$��e�J��)�%����8�cX��Zr	�>!����q���8d�o���#\��vJ� � �������i�
��
������4|���	��\P��݇�#�=��4w�ʈX9�ۨ���N� f���ҞČzXp^���%�u�$Jq�Cj�{�WļW����,�#��b-�L;o*B��)�����+:wi��*�4l���V훪
��Q�?���5�shٸ0�2?.H��t3H�:e(>�-����m#ᤃ�|�j��C҉r�l\������+�������aj�M:'�//�o���r2@���n�?�w�t*N��o|����p�9Fy?w�#;��aj{��C˗�i�K%�ɻ���^�m�M�2���;O���A��SN,��R.�<��[�k�%��	j�"ͧ��rm,�>�x�wM���z���;Ut����x���ˇ}�F����vW��  㮱�m�|�����W)�����A�;�R7��s˗%�ZR�z��J�b<�z0 ��`s�j�r�~� ���&{�%�3��z������z/�1�������>~��2��}&qQ��@�-��%yB�}��T0�'��
AB/�@/�8Jr����McG% +g��Ԗ/��2��V��O�Rfnf8Ȳ�{'A���`ju�����_nT��h]��� �!QGs���}@hml�~���5Y�]Ш{��X�����
?�]�p�*4ar;�O<�R
.'�:���7���GPΎ�(d3�2���/��?��5���c<%��~gߠW|�DR&�-oj��@t�3�� P�+��f�V��>�� ��X�qN�2�S�U��K��deYM��$>�ܯ�r���������&��f�A�mg��۞������aa����Y�[V��(sX^�p��b���&��D��B�5��nmw���;jQ�/�"��7s��g�K�Ԩ���feiyL�]%u�7��d2�����w�fg`PP���53��~��b5�� C�*�-��֬��^ƞH ��c&��B4j�wl�u|�ϲw��g,�[h@�ӐV��tg�Yd8N���=L�������?A��`�S�|0���v���YqB���Ei oD��6�F�Ów��,f���Ć����.�5�L��	QV���}C3�|G.��1`ԙU��'�w�!E:�ل�̞�x��3��B<�-�L� a÷h
�r��u���a������ME=l"��9���~%%�Gt���^0�L,Ԓ�^�0�i1��']��YQ�4AjԈs�B��w�u�����Ծx)�?����0+E�2�8�]0
c�̿E�[��6
�)�|��O(hʅa�/}7Y<6i���U~ �`���ui#6o���o]�}y�V�U����I��C4�Tۣ�1c�+Y�y;�[*e���UC|��E�Zf,)����(�I�/p	@Y�RϮdhye�迹ksr��	o��T����l�Sr�JŞ0\;�P=2��[�?��JA$'8c�%��hj)�U�6m�O�$6 ��6N�0�����tX��}eVQ�)�$TP���cb3�rإ�T�ȦP�6/ߩޡ��Q�a���[��R��'p���o/? �mv1�x�א�쒙}��}�'}��?�;�z9��HM���.��{A�S�T~S$�֭�ޛ�v����Y��Ȱ Vd�,�g�~������ak�(���{�eT�'<��(�<~�]�S7����~�7��Hz�8��5�����x�J����}ߘ�LD//s�	�;����0��,V��D2Xq�%�Q�b]g<6�V�N#��٬v!�i��xk�y�ͤ�WDI�����������8�>��X1k��6�&�r@2����I���~t��4k��=8�xuf���n%��Kq�,��]�*���B~�>�=4�� �;�]�O(d�b�Gw���	�H0�XG��b�<"�6��������s��xq�ַ�͸G�ă���D�W��o!&*�@T�_O��U�d�rN�*LW��=�q �/D�o�)����O�i�ű:!��%�/E"^&i4�y��af+��h�. ���)���VQ�wv�V����(0?��F��,��f��SėHE�Et�4��0WJ��`�5Kяr��$�	�%)��2���g\m�����ɑb`9B9�1\u�W�J�\T��X�/����$�P[m�=9'c1{їM��
�d�Q�+>�Zfk��|d{Ix'%j;�����ЗrKC�~;�~���!� 	&v.�-0&�
�5�v�wwf�c6���0/��#�*�t�_��r��l'��a��𓒓:,����{O?I��Ļ��ڝ�6�u�@�Ҫ܋�ɯ���߼H�;2O�l`���Vؖm%(V�E�gj��<{�y��_�j9�?8cn���Y<��~�ܴ���g�z6�I�,�J�^Q ��9V��NTqߏ*�X�T���.]t���I/�	�znp������Շ7y�9OD
��m%(�ٔY��j��Ĩ�5Y�r$�3����OȽoq&=���}����s6��Fl��!LG��dC�{�$E�����w8W������r��� /��[��K�F�g��ɓ$�P5��w-�yy\mL�kn,�L��f�?��T��.�t~��Crh�+�9mW
��<��
x�-����q-��I����w/!�{v��[��'�ڒ�S���-ws�Y�*нi�m�.h��<V6�n*��Q�p6��)�jISq�mC�	I�4p�TqX��3E׭eA�R@}8�sC/��T���A��S�}c9��*��K�ɇ!�P�[��
3 !0<"�dζC��X1�9����y͊3킏W��
z���_�
#�V�z^'��g�|݈GW�Y'G����Y��XV�'��H$ Sc&ѧ�������n��#]��^���R-��u٧���r�w�k��yQ������Ou�<tw�������?1��+h�*���������Ud�~�T���σc�	X��Kl�)��k���		�6h�O�qw���>x����ly]x�B�&No�&�E�!+����6�I�b��Ǆ����w���z�<Y�-��Lo7��q�u��w��Ь�A۲�d��8X>3�m�-�����fpۥł-�
�Y4ilh�׽$<=����f-%!�$�o�FC%=����@��/W�:��d��&�aV�Փ�_$i�bɷn4g�ށ4���ې���R�	�/d�A8����x��s?����]=O��X�aI�n���(���%N�����w��b�L�۲y5�5�!��sn���v�.Y{�idPH�a���6�F�[�0q>J/��Դ���u�Ј�euV�uٛ-�����䋯S.pn$� �E�f����A���yii�|X
iA�53eZl���Im?�)z�eNQx��\����>���]�ĐO[Azܡ� �؜����\k� ��l���<x�"�1n���.q�>h����7�dD �b��tË��B�5�IO���_�vb��Z��tUX6U��o���� ��`�r[� 4��[��(6-�g�[h�E�UՄ�����N{��5���
]��SGLb5�u����6��֌A���k�9P�B�t��*� ���m�_��mv6)��括Dd��I,�T�����jv�[�����̵s�f^<�l��L`8��h��,윊�E�<��F I��ci�K�J^ ��m�Z�b�[�V�n�x�F�f^R�1Y�����)A�5yߪVi[��£�;K��qChA�,dA�Ky���K�	��BpR�d��Qy���%?����{	$s�����!,m��2�~#V���9���/4p?��p��[*k"�OS��_T�s��J����B��)&������6;x�
�g��
1"Ё��3�W��2o�}���࠺f���0�\��~���X?^)�Q�9��b��
�a@Tnf	^mǭ�P#p�S�b�zR�u����#����A3.�e�8��sy
>�Jl.���6Q�h��D_�T��>��*��T�7���?�Φ��ӟ+���jN\'�J� ��]|�'	���P/�)M2���ZG�T�Ѕ���SM̎� �u�s��uv[�|�>j��L������G&���F��-\c����mոFf�୧4�;���I���|��1;��

�������	�S��������zx̛�h6g���bH��U��#�J��Yz�D�bF^|�"�]�klo<uٽ��5$���um��r�0���x��qwJ��	� if~�"��2�x��o~偛��&���,�y<��er_��:�7J�g�l�<�~l`����\�R��|�
DgG�N�����H@�.�o�G�X�}�`�˰����ueڽ�}~㛔1Q���O�9�y���tf˟P���e��)�9�ϕN�Mr��.�Bʞ��4�Z��^�n�ʬxl8��ɴ#h/%�k����1 ���&�f�#PN�+����xH�8��h��K���`zW��l18R���`9���b��3��ܲ�ƹ�^�W�fR�]�9�BNv=�o�Dt�zf���X Uv����/��2�y�By�~�K+�آ^w|����ϐ��E6K�Ű*�i(�}S�p2��ZP���ZPU�����0c����r�?o�)�ۺ�����Vo�1S�P}�Ěz��7�.�Xr�8Ȱ���_d���	1���n�i��p?7�LH���n��>�`���E2������֙�9����5�v��׏�Ґ#��w��HMW�IfΌù�XN� �,FЄ}��M�aؙj���7��K���r�$��:�~��8�95��d�5U]�uG�#f,�m1��@�`B�h`��CxD��
T�4�����S��Q<�?��U���9��ck��а�;z'@²kt�!�X�����$��1, �@V�pD�����U�\�H�,�*I��pif{E�M�-_�,S��V�5[+�PMM��� �Y���%*���./���t_��45z�è ��95�H���w5�6�xAz=�bHcb6Y����y��_ˇ���}�����n�ϻ�\�RX���1�0"3'3�� }+\'V�Kw$,!� �b̧��j��xstH�k��V�z����-�2d'�L+�Wq=�m.������WsDe{9�ȥY�` Q=U�MWO� F����v~��0֋���Z�A�@�����y? ��p�H�q���<�6>E������C}3#$�[p9�3��2��~��Eb��4���Y��UIs���5��T���zFe����)�w��ʿ�J�h+c:�e�P/�%��?@A`�	�&�k����h���u�:R�H͎�����a���G/�V����m���\�UZ�Z$�l��>�Ж�"i�=��c�@��b��`��AAu%m	�x@��iO�x��dƜ �һ���%n���z<�S��"u#�u�S`���{M�f�OWe,��"�$����[�iR�6�T�`�.��ttl �?��������_��%K֥S�-�e�͚~+�u�w��!�=?>��D7�vX���G��������B>\�`U�$
W��f��laa�����}TES�d=�wG�n!�R[[�T��ƍ[��\�� �a&��8#v�۪�A:ڂ������ΛW/�3�+� �W�pT��,_�#�YPt��HA�\�^_��j��3^o���F�-N��FM��K�L�������~[�����*������-��n��|�7�7����Ш\�k�����E��+嗜��y�ĺ���u�(�o�js�{Z�	u�1��@I/vעa*K��a)��e#>#����)�����#���ɺx�?�uf�&�%���1bAa��ɱypC��[�\���;#�js�7P���q����x��s�}e�N��5�����
H/@ � ���ۧ|i��9�iE?;j�F(L6�獩���9@09_���g����!���P�aQ�%���?I�O�'{����ˌ �OS����T����(!z�T��,�u�[�e�Le���f��$�:v�ח��!os��6��&gh{��&K���A�S�M�|j_82Lʱ�O7j����@�xZ���UNb[��d��E72���������������#����V���� �~x��u{���}��ׅ�6���2�3hH���zb��̥�6�T{4M��YO��q��9�1�E���]�K����( ���͗��-񌠪�	�^�0�^����8#P����S�]�Q����G��ZK�GfFCZh_<�·�p35�_�;�p����6��$A;��fW{�G��5��bc2��۠�	/ Xs*���*�W��7�>���c��V�7}�-'��IL�+#[��������4hT�-씁D
�������\�\]o�ĥ�