��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`ne��kxk�\#�4�b�z���w��+W�]�:�q��Z�U�ۧ�����?���,9������ ѓy�^ϏPg���T����%'>&��,�f��;s`g�q��:2@���6��Wd���jc��1�E�Ǧv��r�n#�@h`Y5o�a\�y'����8$�GCҿ��E��"QJ��Ѿu�����H�Cr�9�!].챩��,%�MB�����1}G{ƿ�7Y��P�|�f���7����!�� >�����ی=�W���-1MGՓX]~c@W�kPA�ig���~��%n�:��`$�H$7je.���>f��?*y
�m�Se���ly��EI�I�ghGPx�/��خP����LC�)�ʲ�X�1�Ƹ/`�:�7B��^[��Ju�l�۲�o
L�ؔ-�d(*zw0���`W3�`m�� f��uI�K�e��k{���쒡-�P��k��I�J��-ʋ�2���x�췐s���t`R� o�N��{��z����}�Q�3��ۭ��k�[ �����6����ӭPcI`@X�2����D��i���q\jaШ-�^N�����L�8������j=�W�<�H)���]OgmUC9R gU=���|N�w��|�l�D�f4�'3j>�eM���w��vIC��^�H��S����*(F��7)V�\���%��w_"���^tw�X�N�����v����=�6�r��'�{���؛<�6z�gE�m�Z�),�EM���r����5#,٠8���Լ�q,zX�3�X<k=�E!�o����tii݆�w��S>��=Z�/���lv��c4�9���X�nՑ`��1I�����\je>�i��4=�M�z��~
�xhK��j��s�K�`��m4����6h�+��ٚ%	BJu�{�����	#�
�h�H� �P4�<&��\�Y����;*P+h��R�Q���{=�.vǔ��������x�V`����<��?&	�n��ZV�j���> �%�,eZ���Ta'7d��Nx��41�����
o቟�6|pmy�K8�j:�"^D#�,�A#*��W%͇ɪ��'IDG���ժ�$�+��i�Z2dYl3f`5IR�W��
YIAF)$i^7b;�Ĥ���EJ���NS��ί/ˌ��x�$Q`f�6R8|��7�#G�"֧NH�2���C���Xt~���;���|��H��c.���b3ҹn�}�:�vWsN�_{�� ��?5�K�N���6C��~d��&G���������[���ӭ�~OmP�!}p-�w�(�����v�`9��H�=c	o�}��#�C�3����3�M���x�#���2���K�Q���z�mI��J\&��G�� !
�!�@�⵸[�c�K%�c��F/��h�G��3@K�wU�&��|,̨��9���Ҥ�H��/?Y�59N�h�	��|�gƧ'�3P��6�c�#ws�2��ޒC����Z�R_/����m��=(�������c�M�v�*B���Gyӌ۳94�j��
R!["a�1�H�"��]r>���j痱���ڰ<�����X�z��QD���V�H���g��f";|=���|�ڭ���ơo�H�Գ���4Üe���n�ġь�y/�[!��r����a� 0�讐��?~�+(V3*����e��@.@L.c��r�l���V|�B-�JMa��l{N����ǫ#+xu*����Z�ߓ&$��r�+�PFv�P������9�Sࡲ)�=�7���	��Az�k>�X�k=��݅��Э�qI"��,z�v�m�nJ�w@�[�\.�w��ؾ����R�( ت�GA��fŝ��R|v`�*�mJ�-}e����.J��������}�������л�t�Y�J��k_p?`n����lH� �{��߼�Ϭ�����\e����g��Bu�g0�s!��:���+O��HT4���]����8� l W�v^�yɬ�'��䠅-�s��e�^=Bd���yzu��5�n�S{ꎶ\��x���Di�\/�����)=������$�(t8S�+m.�]����
_�;m=Yu�ɥfA�y�P`�^}/G�P>/D�qԜ��F��&&���|�B�椟O���g�U��j����H[�26�Y���콋y&Dg2Q����?���K�������6[Ji�U"����~�g�w���*g�\1�����]<�u�w�:�6D�>�D�T<�P?wtt\k�#̎=��k��eqr��h������q�[�oM�l��ݢ�}e}{DO) wܹ��o���6Yw�Q_��4Ըi���7�&�����ZI��Y�ֵ�4�N�,|'pPv��.�A{��-��w�O�]X!K�9AxZ0О���-�!�^[�&ɹ�ə������j�D�Cf���M
��* ��_����7�$�wa�K礢h�NQx�Aj� ��L����t���]��n�~�o�悃�*ز4a1��7�9�e�����+�q!欙�AY��aKI�-Z41ua�S6V�<X��ZUx�9-�8k&o}��v�<~4c�]Tx>.���18�r����Fd{��1�4 �� -��g�v�I<&+~8����M��[������0���C`�fP]f��-����Hx!SGe^�=Q�ƊE��O�P������É��ϯv&V�y�i���C��5Y�Lm���yUs�Y-����뛽�VM�b ���(i@� �~NDA�t��u���wtǟ�1��&��>��5D��闡Z=Tِ�T�Dh9��7������>i���^E]�0+Z����#E�� �A���Hdڈ�;�n= �\I�xjz۹21�5������]��_M����]y��{�����s�v��.�T�_�km�w��=8$"#���;^k�dR���3{p��S�����"ޏmDY!{K��� ?<�`~Р ����ٹo{J�'���:
�J�v���ba�BE
Z��u[���t��=m��Db��?#l�e����+=,DIJ��[ ��2+p��{[���f K�_��L�ӛ�m�����(nj���u�K"0��yɈ�78Ok�]F�h�����4F�,��z�7?t�+4�B�A��+)2��%W�n�#����L*���۾�$;n��Z,���������
.ZG�!�).������Ab���R���k�v����ܛ���_�y���)鯮,X�آr �  �G��]�a���-�/���$�wkX!TW'i(w���ҁUr=�_K̃N����zt\}k����ʱ��n9z�1��Mv��/��ߗ�te˯���JzxM��Ɠ���ɀ}"�����R� �#�
L:����8x���V㸊ov��
Iۋ�+�����Ē< �}"��� iR�e�����t�@1T)���o���� �k�����/zp!wuA��a�eǿ�dld8tnf�j�a.U1k����)kE-�q��]RR���m�0�ssW�	�~��O�� 1U�!���e�:�Q'M�o2X�b�h][e<K�z3sXʗ=[�ai��ѽ� ��Kun��Ҋ�[���`?r�R֢Q�w��I����*�H���)��;N�}����tI�W��Q�#���\K�Ie!�5��B���/J�PQ#EC�ހI��FK��y8F�q����\4��ܖ���9A\�7vװW�����[l<Zn�V��5"���ĳT�(�����?�R�멘4�j�{��"Y���^�����)���ʵ���C"Tv-å��>�nð����h}U��(�#zJ�M���ˈ�Xݖ��3��ih�B�h�cɛ�tF�?$�EtO�T��!Q�58�!��l�0	����"yS�I��Qp�u)	f(���N�B��Z0G.r	�0�\]!i?�Ń�%G�<��uM����+�����P�W~h��Z!�6!��`4t;Ծ�%Is�r8�(%�L'�e�&�)S�$���f�N�G>yS�!怆O-	F��k0v�;P�L�☉�����>���Qs�����ʐ8j]���:��ݎ�GH��01�]Pz|FMA �y="�0�I(U�[����Dcmn�S�2���|;rV�te/����[�PW$K���=z��<������@I��8�F��R͢��Ιi�&e�����B';��#Y|�A��*����37X�� �ϲ���<ya��fT%