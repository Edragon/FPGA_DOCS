library verilog;
use verilog.vl_types.all;
entity exp is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end exp;
