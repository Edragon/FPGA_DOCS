��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n�U���%^2���/�S�r�K$o}(�ī�M�I��)��*T�v�U��LoV�ќ�yk�c.�̂yI*vY�Bo��/fu�����T�F�2&���NC�_�	W؟�6�9��Hw��v��Ǜ��w�]���5�i5�����%t}�b��f�ܧ�θi�|��}��RMgiB��;�J��
(S�q��|�8�L���o'��i�5W��Xy�R�:V�Z��mCИI$�
����ǖ%��w��������,���+UU��]��+�j}�Y,z|�0����K� Ϥ5�Ŧ���6(ёR%���6|�g��#D�L�G����6���ͼ&�G#BN+k-Ğ���a��>Ǎ�V{5{�nXB�Ғ�P���9�K�������g��01ԅ��P;����S�tN�	}��U����+:�ǻy s���Et�=�e��-�)�f��=�|\�6/�},������W�ۡ4���ҵ�{����i��bV�45aܾ�5G�[�_j�;ɲt���.w�ei�Y0�Y�n֛Մ\Qk��hX��}��%^�}��w8XЌ��������Eͬ<��89p&�7��}֓�Z��	��B�08�)pN5d��4����`�w}�����h����rȯ���ŀei�BN�!��'s�xS8�)Ɗ���ʐ�uP0L -���k���wm���Z^�;�ˑ�,^�.*���_�����K$g�_��R��?�Ifo��wU3K�uDi)�x�liN�y����<���`����ͯ~�c�� �\�ި�P0z.��_�P��jM��,s����5���lr�ϟ�^x(�.�~I+���׸4g�g�+n���ީ����f
�<��D8����O,�yђ��p���NK�WA�`Maw@�)���n�Ҿ���v��{�Q�)���t�ʟRFs�I�u�*�m��I�o�{n��?_��_�?3�S˳��Tmﾋ����<��A�A��e8~ܫ��g5a�4��7*Ϝ�e0�o��Ȏ��5�M����x]���9����Eo����W�o6�b����s:]+�E��l�uf���z ��<&�\^���Q��ad��L�h6z3sܶ;#[�|�b*r �c���j2��u��b7��,�O����^K��yL$��h��S�r�*O���Q�aTO4��O[�?N��j��Rg�/Hd3W��y�����z��������J
�0摄���Sp���l�A+d�����CDi|�Y4�u����LV�B�H$��I�y�zu.�!�@�`�=��T���zQּR@�<0��oþ�ÊYܽ}e�����Q�Z�f[�O��ea�آ��p���
��NvG�V:�#��#K5d���#��8uPH��Y�bؔD#l�Gi�����?�H�cׅ$dj�+Lim��m�{g��
܇����h�*�|O�D_j�i�z�+��O�x��{���z�I�o����s�y�ŭ荈3��w6M�	n��*�?��ox�����1kͬ��\���g�{�rOW45�B�y)�|B�,��)���{� �v��;ZN,�� N�R鹼>�4�4b�_D��µ�v`J��0.��$2*�}v+�����+�0�Gi�)�ui���"�RqYP�DS]Us�m� �a����S���x��l���ć�
z���㮫8��"�u�lґ�qIT�$A��Xa� ��[�/O=�6����v��a�؞�rFr_��*VH>�-������	��s��gD���"�$>:8����1��f<g(0}FǕ$2����i�t�p% 51/��&�Y	�[Qo ���WO�䵢��j��SXb�DM��OT��5J]H�ڞs�J����2� �s�*�l�{����ǜ~O1,����{���k4a�N͈{�J�,�ʔ�#p��r}����u;������!f=Z��K-�D�x�Ql�?�7�{6G�H6��M" ϝ�\��;7@�[����pDa�Ͷ�:�ѪL�������[rI0�Jc\�2iG@���\�X8&����!،�[}��r�@�2���ZX�<X��!ul�V�Q4��ve��.���I}zx��3kN� ��w?Ho�>h���u����݈�2>��Y{��X���<e���V|�:U�XG�RhF��%�a}A�Vd����Ӥ_�%6�,�VF�];��{�D�X�P*�U�C�C�g�{��|:\�I�&ۓ؆�=��0|_����8�����
PW��rsvlo�j�i�؅�ʓ�Q.3�6�z��C�:*���C>�B�(C:��� ��]]{'XBVNLþ���t����J����]J�aIz��M�(�&<١��m��m�]�+����h|�a�e�!��_�O�j�����J��7��i�,�:�?w���G"-�T���-h� ¼V�^#���*-Am�  �Y��eA�I�z�>��w� F�8`|2����y�:*G��!����ń�����9�w���25�����q̙#b��؊a\�|k\Q��Ґ�"�\���!Bj��!+�%�̸��5F�-
�,�����6{�D��W)wgV �gy�~�����[��ߗ��?G'��8��i�WE_d
(Uk��F8�R�YY����Wȧk��JG^��ʀ0��ő��iP
Iж9��.�T(�P�����l�jC����|a6�V��O	A��v
�S	j���r̮�] `VXJ�S��)����	Еy��<�C�/�G�TY1�V�'��+ώ��8��g���x*.�	�e�Z�ל:)�����Ɣ��:��4�d��G��p�f���|�s�@���<�щQXr���_�Z��B�'�1�]U��ɫP�f��j��D���d�X���b��^q<��D���Hs��'��Z9�Q��Z�Q��6�;},SmL��i��.đ�H'��D�7գ�ƅyȋȄbm�e���ρ�� �ٺ��|d����69�ǻu�q��;�!�֌��>Gjn����\B��XM������k��a�
�2�C-vT+L�ϰ�V��SᮁsDVU���.]V���.���,X�Jȿ��͟�k0ם��� �p�"��P�b2��׿/������}e������2����a�(�����wg������1�Q�0[\��R�FX(���4�o.lΆm�%��J�lƖ��֋�";��O�?���*%��~�hd@�	��6f���tqvt���d��dg��6{���)'���d\���|Bf+��E�Y"�D��=R���薒�O1�lͣ�z9��TD��l~�r���|�&&��󟜪�����e�'*2�U�"�Q�r%@��ёIӀ0�ř ;?��Oy��c�}��+Ǝъ4�?𣩐qv{�v��5��B�s��eNv�e�e�$��4\��`Ô��T�O�vw� %פ4���h�H��.�tJf�3�漝�k���!;���m&
a��j[)�h��n�'8nF&y����-�Lrd�U��*q&"�dߵ�����.�G
�{
��0m��L��
��CdSПT�M+0�ģ�R=X/�`r�q>����5�� r3��a�6Y��8-�Н�T���81�-��Yp����;I�w����uHp	n�\�=�CH�n�����L�.�#B�gj�
���Ș�؊�wÝ��dC�4�����%$סɘb���,2���5mUU��M�"4�j�ߏ8t[	-C|ת�I�R��?]h�����lH}����2*Rԡ��x-J����Q6�G��z�#�L�ɔ�������U�Y4�7�oݒ
7���W\��%���9�&���;�8U6N88�}��qF�����֓#s�;�ve>Tw��35:״Iy�1��d�� -�8N���4��b�l}n���,������5l
��5�qH�����^���pg�s���B�0�:q��^f���3򸠓!Y�"����{������;+#�3͏��<��q�B����1����P_��j\,���8(�{@�]&�#�@��N�B�f�]�Ҡ��~���؛�x�B��hПN�x�� ͬ�(ܦ��_���r�:�D\������1�>��E�o���74-T�;��&�d+If�;$.$���E%��j���RL9N���pT��^�K�|�=t?K3�(O��u�hϯރ�v�鎶���L����ϕpmAE�}��ĘR} σS�����&^,�����l��XP�Ι��2�����'ڰ��g�.�GU,~Ӿ�D,j����;绠���l|��z�Ή�n��Y#��]��Z
����=E��|Y����Z`�����)�t�~�)�E����e�5C3)[K,�[��:�W��C�O�fn��_	���w��5�8���N^�5r~�bs�U%,�1�6����RQq����)s�U3ZI�Z��8$�����+E�+�z���Y�-
��/�<>���	"��5(%�Ǵ���b,_(y�[՞GG�| �A$��9,a{�� ��W#e�Ig�cO��.Gf�G�e;���3�]&!�Ʌ�;�-��)�Y��`�Gm�le�Fd_�)j�zʸ�Wɷ�6(�PY)�]X�W�"�PrgS�P���V�d�I�Ix�
c�sB�191�Gn�\��x)�A3���!D˷�Q4_G��I@h�n�z��Ԡ9��� �'j�g�)j:�C�m� ���=8����ʉ����w����I
G��,Mڨ�L	S�o�~���T��瞆sp�,�T��=���Y|�nfo��+;�w��u�F]�����#� 5��2,h��E'W��^�ܵ���P����Τ�<���aC%��V��ֶ<\���"��P\�ˤ�o����;;v*��0�)�#����7%�zUP��W�)^�X������&V������2��c��D*Ӝ����\�&��d�EHXGg�8-w,�Z�?b�
	 c�AMJ����D�2�9,�8�@H�������Z+��T����^ˮv���Ӿ�_
Pڑ��Ծ5��;���e�s/o���}�>UkC�U1�g��B�6P������<�K!
	,F���&UӀ�G��E!�&����7������Z�h-S~YrA�qW���E��%fz<3�u�X7�B��@$�@A��t8��a��*�JV�~����|I|��u]��{3=V���Ϡ�F���5`�/�d�qr��-mgme��l�]7f85�e����Ф�k�2d(��<#�v9)?k��@������'5���q�$����3�_\qcq~�u�^V�$Ytv��Iƛ������5,�w:_���G,Ψj��<i���ut������.����Į��'��l���t�� :�ʝI�l����&�'F�7�Q��Mx}�K6�����# ��j+q�Ó��Q�:�j��	2׀_����K�K�}l+�g&�Z�9��J�y�sP5�%�[8QB:ۆ'H2]L"�]��øǆ�}��Z[�=*��@�<d
@��Ѣ�?���#ٵL��E���3�/7$p�i����{�	:�$*��U�@�\5�V*�����fm�]c�]�d�k.'ِͬ��� 4���}�2�:��IR��OG.s�آ�3�C���!�7 �Z12�������L��ܿlٛ�
��-=���n�m��G�]&к�+�H�0��JFgn�N�������r��)�u��-�7W�:�X��m{����-�{�|Xo7�r�_"�ѐ\�1U�A��қ��"bȗ݆a����)���+�����J;3*��^vc��n��} ��Z�d:�"�6�t�m���D�O8�a&�"E����'D�ȸ%h8��׋����Y#�~ߌ�5��E�f�(�M��2�[i��������V|����I-w����/2����-��i������7��@�+��H+���&�+����o�^�b���w���Z�K�ysj��ѯw��}ƭb��������j�F��Uv1�~�q�,@��z��g�`٣���C}iq2SA�Ɂ4�?05��^67�� ��W���фIN���Z��_�����D��ޞm���G��'�Z��j��F'|���d�H)5䄥S��׈6<'�3�Bk�4�NEx������H�[���n���[�ځ;�j_���|�@:F�Ć�zR>���`�0Itms�v���*�5	C�~(Zj��X}��^%%ɉeÛta7���$x����N�%��]Ƒ��WMŚa;��h��0Yf�n@�_4{r�(��3)LS��(����f�	�rǞS\����e����䊑%���U���L��@g���n~�x:\�R���+ɀ�]����g	�i��Q�ˡ(�f��}�@�Š��v���n$aԴqk�О5*�Gsv����s�Pf�A�D
T
X��V2�!z�:���sšl�<1�,� N�2��6��T�GA����k�tֆ*H`.�g&��#�6�_gM`��k��V�׸3�+y�m8-P����Ouz���ABP+7���隢���c�K�,��y l�k� �H���z�������o�z�g�c��U�cN_��΀��<�"�6Q�#�K���p�VQ���d�-�9�TX������j�0�?�y�dk�}bi��u?�c�w��'O��nf4{��0�1<�j\X"�݋��ɜ����������N�k�R�8�F?C��J;��.\{'�=���KӒs�Ϲ�/�㵾���[��΁�
F��N���=�q?f8j����÷5�\�v}�I�/��*��iH��zi�' �Aq�b�S�4�4^�7�����,[����V��mv���C_�8W8�N�f��4)��Q�>�{�ԯ�+�.�)��(�q��Cc;��I$��&�N�	L0� ������洐����l��.+_\�>^���`�,��G�Sʈ������A��|7	�'��5L�����et_��?�|�t�7���qZo�|n�ۀ��3^Y/��(�0}cV��B�� �t3�F4�X��X1u�Z�L�T<3���Օފ�Vȵ��󊶛�6��(��RjY�Y��U'1�5���_e�B�a��
�g���x��5t��ĉ����X��r��Z�u9[�o@A����� c��]���y����l$��u��xJKG�k�%�
}��Q���l���w[��&�0RZx�V5_����1����*_�l���Kl���Ao��/S�f�y�w�鴺����T�`�Tk�q`�\tI�8�� ࠭���ϓ]��7x�g)A4,�8�Fu�>5��������u��|���a�����]�6�5\炡"�8A���p�8��S�W�w�v6R����0޲ �qy�
���8/K��0% ��i
kR��Y�Н��s8$��*�e��ǣG��#؈�?M*/8}h�N�f0MM��u/R��Lp�M9�
~��m27����=��i侧�QG���{i��J eOCo���'<�2��&p& o�eN6��4_� �G#KK�R��3bR�{3�m�0 _Z��(LV�����k�l>�q�W����B�j�1�}!rp�"YT؜���� ����+n"E��<�x�.�,�ȋ)6��٢l[����gU.�z-q��_�ҧ譅Ɂ��� ������
F�l¤�]��yH�^�^= �
%�x� ��Ջ�O�aH���8�_��7{�}�#�����/Ϥ���;�i�h�+�Z�L����`,������'�!U�?���r()���{�ci�>�?��F��r��a-b���˛ ���>r�a�-�Q�2Z��A0�!¥���1=����F99�$tW����@���y�V-���ʁm��[�s�͹��c�I�s}�B,����V[Z��E��F�L��HJkW������NX�R-�-!�&���Hv�Uw@M�ך�d:R;:i}������d<��]�;���7Y���ׇ�$�}8P��h�͛�y/�����M��U�Gӕ,hUa7�r����=2��A����S1� \m���,����n� W�S�S�W�ԃ���O�N�4�R��R�ٱ���,�R,��	���bT��V���� O��^��͹=I��FM<�s�.��Eu}��7�kl>���[O:2Q>���GyUX�����v6��1��A��ī���h��cڂ@�aa�I�~77M��c�v�{��h���ʔ�v�(���*׽�̸nΗ�����^1�@)�}`R�RGe�n�_�^�d��w�vm*��	4�&�o<]HK[w��rV���۶m?+O" �HK�G"@D�e�1Y'��T�V��]��U"�h0{=�=�3�FHd�>d�?:k��3�J��e��E�?G=�7��͵\�,�<1�dن�iJQ�O�H	y��Op�Ã�,ńD�vH�����ua�2�$�A��Y���Оx���.��1��aU����ڷc�p����D���}�T�7��W�T��Q��͂m`���[1��ak�Z�vdK�+�'0'�d�ɠ�Dk��p��KY�m�C!�$�л&�LB�;�[���e�v�Cm���C+�(�j������'9���-��9��'���d¸��4tCoS3�@���H�Zģ���4Ѐȋ���*Z�t���cKLa� �6VB}Λ��{w���l7����'�K�(Riga���$s���ơA��S��⧩"���Ե�M'�<�dd�*V}m�vM���j6�)N/�U�� ��~������U��a"�7#�FS���Pd����$�G����)�w����E!��0̶j+J��fZ��y8J6X��ޠ_;��38��DD��#��c-P�������	N4��sc� ���p�}�����H�~U}v����ㅩ�Fr��VP7�SF%JK�=[ ˱h��fR('!f0��Ҡ�&S�L�>K��=f�\=<zR�U��Xچ���FQ��ZF)�����b��CZ��t(�@�K�'O���9��٢��.�\�Qiu���"�)�*�/{͓^�^(�Uw?�>w��>��a���4m������7��wg2!�w3N�O� �6�i�V��s3�:�+���4ʘز� �� �����D����Pn|��L߇�Q&��+�6�C]e�S�6,�g6$e�n-po�l��ڄ=���U���`���{��͠	�����n;���w�uRୁ5�`�=�Ǿx�
	u�mw��m?d�:�jrb���|jC[e�#nJ:H�Y��a���	w?�e9����Oӿxp#�fT0Y�n��8V�@N��%���S����s���qc�Y��%w�p0������Y?/�x_
��X49���m� 42�;�W�*��;�#��0챎vv<^ȵ�%I�{fZ���ۄD�52��@�KM9k��ᱢw��� ʞ��>z�)Y��/Ͽg,��	��CDu��ՂH'����9*���ݩ/y5ߪD���
�H)�c�:�'@R�����i��B��)(�D>��"�v��+`=���n��Oo��,9�O>�f�YFȊ���5LF���uޠ�ItbP�Lэ\��ĔVwyʱ�f�"i����xZ�ՆK�W¦�`�����y��b��h�ta6ט�ğ�Y��Xz�}W>e�E����<l9�6ɨ��2<����U��,Д�P�'��X���Ρ�����,ĩ�
�[��P�}�ePf���7��鳧�b�֑��
�[��5�i�Ce�1�iv7����S�d����|$��X��N#O;-RT�x�|ޢ_��� O�H��VB�1��A���)H�I�\��m�G&H�_\��Fp���`���B�����wՁ����>E�s+�g��f5�}"�D�di�׶�ƹ�S����7g�P�z6�'c�����y)q���)�>�W�)�����`���FE	�p��6D���
�`��dʄ�ҁϟL����)8s�x@n)D�O��rJ1�k���+{��x���0q�w���� 0b��$�}�-�K+h�I�	w�[���T��m�n�U��g�σ4����Ҵ��-wY�_��(}j������_,��l���!�3*��������2�Xo�sX=]�N���� ���U+t��9�)]��D�ۗ�-o���ڄeϾP���/:uzm����_��8Gnjɖe7<D����!���:6@K�p����1'Χo~e��n��ǚ$|�Qi[����v�\4��Nb<��>wxG���K"�i�m�C���ٜ�\����\��X
�&�ۓj��`��3o���ž�I\���á4{w�q����A���S��`�7���0Ԭg���9NS�zJ{hʇ����5�\P������o۳��5ɎJOmś��E�Ղ�6�x�IϪ���� �R��#zO0��s��@k�ńN���ɳM6s#ᮩ|oGxg����N
R��	s���y)(ky�(�S���>�V���3b@�6�a�d!�wl�}3��z��0�l�7�~ ���e��g�>=�\�Qv���`B�m���JJ�V�g�q�	�N�&�1���:�D`9�fs���k����U���O����b�܎�\̊�3ЊG�5���a�g�E����̵��>MqD��]PV�n���ķ
���*N�a��)�Z�>ppM�
&�z!qU�aL��_����!dɍ�
\\��[�3�;�I����J�~쬽²#3B�7���dȅ���XRRr�κ"Ad�낽.��&��m�3f���;��MK�����C�-H��k\���b��l���+3b���{g=��VDxW.�,?���*(���'�!�m�ޞ�5����kIK�V����GT�bF��g���&8���swD8^p��`Yq�}W�-E��&*D
Rs��ϛ����r4a��j@��2�
=�.ӌ��&�)g2b2�l=)���S�iB����6q�Eј��=sǆE:1�k>��On����P�Xx_�#�w�:�z�d�R൨H�� �{��A����.i7M��mh�fS�MA�çtf�!�/+R�{]�9�L/;�|n���q�.�����4h��FB�
t�"��Qӓ�<��3����)�=^;�t��c*�PR�P����:��7*�s�e���i�g(�q��Z�o���[���^K�rY2b��Z)���.g<�:E��;�ݩ��H�ۏ�X��o��f]��0膢������ w����~'_
�[�e	�xiv���'�D��h/�*���w~�-t�(C�M7�2�[�y-a�7��u� L����M������m�̍���.��(��Q�>�d^�г3gp���[X��3�&]*f=5����=�������
�M�)�<�"��jM�Ԓ'3�%-r�B��#lb	$ %���SS�M	���1	.�̗��2�Vʸ��D��+V�'�,i��I�'� =�VW�"���(�Q���c���~D	�>w����J��X��?s_Q=�U>�>{vC˻�����D�k")�|�!�l�K$JrN�����ƲI��r�T;:֜k����D�F����)�����ogh�W�BC%-Ii_�(��i�2�Wk�a��jG9���ݡ�\����즻��u|��l��6�w�2:el�]�`��JB0rQ��۴1Rp���&<Q,η��e���mhQ��>�D	��������԰�p`�P'<�2�zV�iuӕ��L�vp?�A�a �R<�x+����x]��hh�t�2��-4�0F�����_(��s�@��1Rv{y(���\Pq��>R�s�q��Cb�}�hq�IV}�X`�^2Iȯ��	j	���g��_�q�^�ډ�����^� �0�b���˴���E_4����`�x���v߰w�{m���a�yLj�DB���x�7�[o�*����*D��H_=�T�#��v�/�q��\��ꤞ/�Q���q�_������d����*e��[�\��.�	�厧"Ř'�f(�~�؈L>���P9-��S`��e������a� Z���T�/����vI&Z�Rmy�����M���;H��)�f�C.�|�xFOl�v���yfc��W��2}D�.�������p(�O��q���0`�O5��jd�S���M�I���\���l���v�����i04�/�s
�X�Wen�5�E):dk	�3J��1D={��-�l9�x�wF����ᄢ����SH�Ȫ�=_��u��NZ|��_M�`j�	uc��2��8t�zV��'�f[��Wq&Mʧ�~#�K�
d�W�(�zCZ����U��ဧ.(�{=\�Q3M���2��!���U�Y|w��`!T�?�T�FIOb2Y���D@[8������?m��h&�dЋ}p�����P;�w���,.d!�T�6�_n��A	j<w�U�F���m�*�w15E�a���br�cE:ǋ�O*x�.N�Y��:]	7]4��g�ͅz���� f�����RsR�{|Z�]wZ�p�n4�@r�Q_�Q�2(�zD<,Y���&+����%*�3(jR���W,*1z�#�OM�>B��wp��n�g��F\)i��b�͏�_��
�ﳛ1�h�r�W�p��ec�G0�Y����	[��&��gy2Ryf.�d��4��Ҙ�����Re��o�cB��gH�X�qV��8t�5Κm��]�ORbl}:ܿsT�~t���Jf ݠ��@��T�G�[Sq*�̌[�!@��"n=��0�4�栢�Tr���>ސ�S
�V�	T�f��3anyc�O)卤�`��7%���mA7$�,�.e]�	����c2J��U����/��
��dq�9;�ɍ�f��ǭ�˂�L�ʻI��S�'�e5��'+�����_���L�t�H*|(�;�9 �@	���|�b#sMD��ocAh��ς���Z���3�}�Uc)F%�Ryʵ��l�N7�5ɖ,�V��潕�Ҍ!��PEj"-(����>^�"� �@N.�x�CF��ٰ49,mjx
��y7�W�=%�Y���=J	׋v�T�]�Q��z�Wr�`\��CKf���i���d��h������,�SB �g����_5� 0��Y��*��$K�!�xe۲xv��e�7?쩎��IY0iD�bI����jO�����B	�X&�:�����n�7`��4�;_Oj��9.�}�R��j�'a�L#�,r�2�ua�褆�X�{�.o-��N�s����QE�MH"�vI�$���P��9Bc�z,EJ�>���+P�B<��1/�4T���d���a�R�lE���\fTg\�]K�mfd��ک���}�e�� 3��]:�ڤ�ܼN���$p!PT�Q}��zC�I�0�a�_6�\ev�T�	@s�G?[�>��y�6����^Ϧv�j����'���!�g��j��d�ݰ�W��%�&���T���`�6�e��i�_��f!�U)b��e�����~�%vFB:�+�����5�񐖮�r(�R�A��cں-}ʈ]㔟gl"i�r�g�=��� ·���9Ў2.��T�4�f�����ޫ�R���&aY�z��߷8jŽ6X�)� �Uk���#b���g-	fF館��{�����۪��fZ���M%?��g�~���3���E��ҔA��:�#+�>Z�G��ް����Y��փ#)I`~�c���X��xiU���"ܠC/@�L � ��ĲSﮘf@E�5�k���a�5��S6�`�U��+�ߗ�S������R�XG0����ܔ���Ռ?:���ԣ���e���<5ǫ4i��"JSi� �UW�B쯝F���n��C��7�O�i�y`�Ƭr�`,��y���+����ͻ���n�W�[&��m�-����&� �ѭ{� Y�QѢ�Ȇ�����N0~r5(��aъ��]�1��~KUR�;B
^���
[(�1n࿵�Z8���{Gm��o��
��6|�f�UY�-A�s�>�ƛ6��J� ��4��i�Ģ�L�.���SZ�W^}!j�:�jP��N��a��A$�? x�	��S�J�����5��@ �=3���0 tp�-���a�K��ݬg�rKwDxI�$������f��2����ڰ����v�	�����_�9���)fq�|�������{C,�� GЊcܱ@�k�m8`����x_R�n��V���?i����K"��¸jl7w�"S�`�z�{��^8Ͳޮ�o"�!��s�*�L�GXH7.rO���+�!(c�
|'�YF�xFW��fˀ9� �U���F���nHMWz�����6%w��ڻܿ��[HTܔ���Q����v��ʋ�<�^�E��|bQ1���	<�w �E�oU�.�p�o9�\��gܟ�ΝQ<���(-h#[AO�J�	�ͪ�}���^ޞ�J2���U�}ƭ�(7d�R�d��ڕe�5R������_'�W����H�h��b":��!�a�%��/H
I/-�@��i:_�{�v2�2�������S���и��/A�@IFH�8'������ڨ���ޜ>��oG@neR#�:�ߜ�á�Ɂ��M3N��V!j+SzHX'7H���O�#!fҽ�ajK*p�w�:H���J8h*�_IW�冕��q�g �G�˾BH��KU�J[b�6��T��VIM����J!��W�\�S�H)1^�Ih����@i���Z�w�\S��q��a��B���0��fv	�荝� :���}�í��(��?�OD;3o�@r�_|A(��͛�`+���	 ��aq:\�:�Z�[��B���=Lt�#�ɨ	�78�ka�4-$\���'0߸�[z�,2���ži�� ���{���`�pU-�.Hk�(�
��i�>3o��h]{j��i��+�<9TS9Δs��o�$��E���$S��6�}�B���zz��\�Ŝn$34�Ub���:���
��I��@������"��S�ʃRS�LN�݊��_�5���MȳA�SR�A=_8������|�l�IFm}�N
2@ʜ�]po%abekL�����N"���(x�x�F�V��A��<j�nc*U5�G��C���a��`��{�l��& Wh�O�B��m��������mx�ۈr�\�腱��TM���Ử:ġ"�3�������A�v��𱑀�c��#�p26���``���Z�G��W�z���7ľ�!���@'1�8Q��E�o�T� �����'�>�Xm�}h_g���-8�������AscQ�T��_����~��m���wt��>�{秞�Y��-�ZV\�s<���?���`����Rq"W���'�]Ŕ��/����+T�@�_Y���K�J�����g0�ý�|��b������j^���H1n芮h�vm�twį�&N����~9�X�Q��M~�����p%ƚ�j�[f���mAۖo�Rk���e�¾�Q��@q͈�ك'=7$H�f�Zc��N{�XoV9j �l�ʹ�D�
�J-Y� /m�l�����jn�0 &s�Q�)��h�>a���)CFzpLN�T���k:Y;��zK�E�oc���Ď��.�/\�����A���<�/�c9�Q�2Ƞ[⿽e�˗+�SuN�/N��c7W�����ز���eT%��N��i� ��C�jrMr����)v�vuj���>�k�s�GhnZ����%R�/Ȥ��3������+vPՑ�c����Ƭ��lY�W�:���}�?�<�'e�,ԫ���w`=�� �9o[�M}��8�J��S�E���`H=�?�+�t��".�_���G��w-iWpā�Ewz�v"�f)<���بO� ����-L^��lȅU���EO��	v�� �;F���Ny�+n_?���t��%��Ʃ��F�A�I`l��2�M�D�u@�7�/W��t8��}����kC�d���)G�4���2�ܮfU�A�8V�EZ���,�A�Vx�)�e��ΒkܿȀ?@��A����a��B
�S������	�!p�n��N����R���un,`����Ia$������e�C�ڕ�)�?�V�-������f������T�S\y��`.�7?���D4�WO�aՓO�U��ir)��҅��8�CȺ��1֬W?6�r�� ��~���`)���L �WqDMG�m�/ 5$=?�QS�4M�wplV���L��+�*�w*�'�]U�(�kw3O%��N���g�?��n�7��V�%V�T�4��j�v�lO�Fg:�C��F;������ǣ����ܿV�}��2�S�X�M7��R�T`*��>�*�U5�{s��=����J� ��#�Cd�=�c����W���D�z�f�]P����=���>l�3�p���m�k�Tz���N;�I�я&I�H���U�?���$�~h<1x'5*�=ub�:_Q�#�SkÌ���(,#��S�[-�x[���� =��lU��.����sMV�b�#H�$\�؍�t����?d�D���rY��A����ھx
�8PvL�:eYG�	��OU��f9(F����
x��H[�W�w��%���	�W�6<W��b��4����&�¬Zх�(m&O��`��%Z���[����M���YW�!���HH�2wz���{:��GoL#[�}^��4���Y^��ʱ����WhÃ�w���]�׆G�G���z;Q�pdRO����1�N�v��Q��i�E�����`+J��cOT��_��i\�e(���>&�Y�S�qg��<��d$�vc��4rE�d��ש�S<&�ö��kT�v��Q�[rq27��7#�TGx=���S�p��4bD_(�HW�J�i	��0����1�f�@��(B��IH��� ] hU��I7I�P����|j�%��.R*��]i��Fz�>�P˘$,�f�qm��(���kmSm�����O-Y~8E)#H�[�u�x��_Y�9�y�4��Xh���P
�l��ȃ�:x���e!��&m��$��aE�2T)�3����#��  ��ǚ=7�< ����GthK)��ǚ�I҂)���x��V�G��"������G̕`�)�����u��DI�aۮ-b�,65����|c���V���"(ۗP�ْ6[��n=���'�R���8I��+f�TE�81k�eX"qnH$5�Ss/օ�8 �H�*�u�� Q�/붺�Y�O�oBP{,�g��9-�G��N���u��\X��Ů����U�j=�z���SzTo3�]3n�9�V�VI�ɗB|v�x��$�T:r>�	~�/�2/UQ����O�"���}�Ed�?��)���hC�4A۝���@�FDg���oq�T��/�����Z~h�	$!oH�q�2�Km�ƹː�X������
3C��65�(���Kۡ�)}�$k�W�'	�Uo�`�%1��>4��<@�a3�� ��c�0Ds��(��I� I��!Vi�H�z�58��Z#�H�DWa�+���C����J�(ߌd*8aKk�uL��#F�aB샂u텺�;�w��-fk�Ŗ�a��ȃ���e��k<���*D�q�w�Щ\v��	)ҥ��d*5��Q����"�1?.�F�t�bfF��%�:�s�.��`0����\%�q�R�;�l�w0��F#�t.���Oӑ��/��A���Uo�q����R��ħ}4s �u����0m�1g��'E�����ګ:�1��p�I^��DAm>�Yܴ�����P��^pԤ��6
m��Uy�.�������t;�R��Xڥ�]Q���[gdVݴ�T�i\�r73:8�E�Xɹ7�b�``/D'��E+L=2�'��ZD_�O��c8Z��a��$*���R;�1n���J�l�"/��/�p�԰��Z���+�T�W�Zw��̾Tp��Y�W��� r�h	E90��#�;OÉ~JཟI����W4�dW���+�Mw�_k$�~ s:���a5�Cz��p[��݃����<.N'���J�Z����"~�FH�H�Z��p{��(������n��3.s7���0�G/�O.�R��|��ղ�/�4���dú���0܊%�wLG3 R��W���>Ǽ��(�qo|�@���.�B&��Lm�ē8!P�,۪�Jy��sK1�*��&��:X�s1r���p���� l媯�ѫ�����u��ʶ�W��kV�Ľt=�ڳץr]�eF��AߚI�h�ݢ����ұK�X�NN�i�|��� ����Z8{�eװO�O�����ǯ����D�@�%W��4]Ϭ�
�!22K{˴t&<�"7.��v�8x�����bO���g=�gZv��#�gBd���y\뜃h+e�M��Iȗ��Q��\��B�O���H%*�p��R@��D"ma�������v�:�tG���~XY�U��f%k�k�{3\Gp6x�U���le)�?|	e�<@�	_��
��;�:���C�u`��G�)��Й��Qi��\��|���K���X6�w����Q
�0b���i��hK����
G ����cO�8���)�w�B��(q��g�V5e�����i�E�����3�I�i�!صa}Hl��T4n?�X��db�f�"���&zl�E�c����+�����Ҫ7�`�Mj�H�w��Y��}6^���Y;g��4���/o�i�y�ˎt"�Q��m&D�P���n�	��[~�]�cd�����6OL�_��l�xY�R��̱�2�"#�>��O������#�*1CIߘ�=�$}���&�8��Xd��єw�cin�HEm ���/8ak��?lb�#n1ޣ'a�f�l��҆wq�T�B�ǃs�@C�Dr����At$��fT���5ʸ�PUG�=�-e8{y
&T�?:�F�}:�}O�Q����:�=��aDqH���g�%��lm*�i����$��'�\xM��.u�~"E�#F{�;�SA�]w߉s��7^
��gb��M�\�ts;X����
<�(o�B�lߚ�v��.V21$N��Α��z���@�i�1�Gg)�*a�>aʉ�v����k'����Jq�]��깍8�*Z�]���ܦ8�SL����R�a=�U+��Z��&���i	7PHԄc��C���;�]��e
��WiZ�K��;4&��x�1]b�f[#��j�M���֚�Ol�0P97�F�f��,y�_� �Ct�C�A�A5��?��@�K<�����
���ټ��)T.���n�è�7w�P�\�F��r����(>�O�O?��,����'L�w7/�S��#�����2�����Пn�tOF�9/|��o����
a�^ s
$7��E)I�� k�\��&��nٮf(�K؆����g�i����R_
N�T���_��E��T5��߆��W�_� ���D6�E�7���Zf�%�1�r�e�!���c���)�
2`�D3��g�B���)E�VEI��3�] ����V�:��Ι���i��F����3�Tw'�GU�4.JMt�K�o:�m�,p2T��tZԺ�Jī!1)���`X��rE���'+�O��-pNYc��L��3��վn��e���KD�j�2���k�ٔ�¤�N��+�v=k�nŅ���@V����}�j���� >��B+�`��<#PШ2����p^ؾ��BUe -T�\��?�I${�xJ[��:�D���ĭ�82=�.�W	g5p����4r� � ��芎!q�-c6�1"�*���ٻs�QG�u����=���AzX�*�1���$����v� Hv�%v�r�L�wRF4g��PX�3��@��e|A>����,��Dn�$�����n �8��������AW�l-"�4eV���N�~�^���s�ȏ�]>g�k�c��$�@*����ʶA7CI.��kO�|���(ͼ�����{���v��"��Pv��8SC*&�D-���$�	�������<�!d���=��%����,(o�T;Z���i������>��H��YB1��2�=-�=�n�qw��J�Fh��m5�	��&U$��)���v(�^E3x��*��#F��\+7���Ri�/)	7�@a�s!\&�8s��_B���p<;F���i8��i����gq`Z4P	C<��2�����F��cI���"��}�&�R*,����C2T��#TO9ы��F�:�����\F(2�s��k�.��Z�*�Ǔ��a�"�^��-�ȷ���A!�5���jd�q�XS/t�[犞i�����ڹ�n��ۙ�]�=ۍB6���,hE���u{���>�ͫEi��{���3�;U�(����g�������43��sd34��ڎ l�Iׂ�5>d�v�ȍ
��b�"mk����H6�6�o��S햎i]w4]봢 Q����nG�%
�}^<����_��;���`nz�T�#��u�']���!�B��h,�~df���8*	۝[X��]t���&�XX>sf��;Ӵxd����������(e��āl��>�9��}�G�5#g7s��z����z��h��-B6H�q8��g�	_,UP�d����hh����O�����6Y�;����**`
����ˬa\^��,����#r�k���!f�x��XE��w�4�Kv�CSk+.����/l���D��z=s��c���;����� �e���'d����k@Z2�Y�T:��ij���YwY��ǘ�\�������-��cx�R�u��N�#�7^��Ѫ��<nѸ����\kt#C��:堽y�m�~}f�w�g�t�C����< H�^��k�$��u8�*c�#�yeLL�����K���4��A��$�?�+R�w��T�ȂK��W���/\O �\��v\�p!��~ybG��	 �xw�E�-��ֹ�C����C�ޛy��j?�O�ʆHF]��U���0$نzF
&AHc��}���h�dd��9L��j Lˌ���K�12ҁ�5$0�.�n+I�2�	Ϩe}f)^���$��"����}-V�\T��BX��A����,J{-��|�K�[��lt�d�U�0(��)h�EH{ӊi���.��}"�z��c�R��H`��?��',d�R��~�yw(��*�����v�WPHf�)�M���#�@�iEv��{i誜\_AU�Ǹ��� ��td�(��ꩦM��uc�W��dVx?�n"�d�l�>��܃;t�/��#]n<h�����j+�rڌ�����[Zޤ�vu����D��G�l���i���U"�"c�s�"�=��x!�����q�g�G��](#�����4̻�
�$Rc�oߔ�і��{?�����S��{;zg?(Y}w����XaQ[���\hꚈ��n���?��W牥��ʩ�0N{�V�yQ֭Yk�!]s�`ʍ��ն���[���5��bY�09Vo�"��F�F��ގr4���~�5�f��ʯ=��^��F�)�����#<�'t���CW{�M�8��!��{~�����lQ!���GC��1����NQ�O�� nZ�i��>��C�d�w���z�L7�K�����"|�$Z��9)
���b��x�U���u���_�l���g���p��X��|�b�ӂ��`��`��U�o���mxӮ����ΰ.^�P�ҳ�=�����&��N�wGi8{�E9�k��'�m��73�UGL���4W�g7��)K�9P����9V�*o�zys�o���Q�F;(������FͶ��=<Y�ؚ�CK,yMy��)L�|���9~�g���N��>�؜�*�\���N��(\�o�ڴ���w3^7s�b�zk�Tyc{����S�
f��9ԍ%�
#��E���]�W/kn~^4%��h�
s�0y1S���Oh)�ٞ#�e��Z��f�k��z(�����S�p�	�EN��=���!-@5��g�X���@������*u|Rb[T�g�G�F�Ex�Z���j�"b;�٫��ԩ�!�.a��56$�i5�^I�n�L���~?��1{q�]�u��wB[��"G]�8!(�J7�b2��&�Gf�q^a��k�"π��u7��<ƉJ_:�`Z��{T�Fx��h�>Ыx���=m����(��Nv��<H\���%�T��R��D�w�;��W� ��ߎ�C�yZ�����`����B�ą\�_����ұ>�]|�J�F#��Z��:� �x�P/%��x��c���c%xC�䤗����m�� �@�KQ��MDB��n����*[ܩͲ��?4t8��:mR�-��!}q�l��x��S�|�1�H�{��&�bQ�^7
�7\�d�q����M�4Z���ª����(, �����S=���UM2@
bڋј/+~��������WR�M��sT��Z3QobMX�)5N�醿q�`Ѥ,[)������@�6r�hU�l�J������V7�3^J%������!$L��\�K/t��YY*=W�ۢ�vW����'O�,yo�(��e���JV���QsBe�!}�\�8?�d���0j��E� �V]��'Hx��*U̺�+}�tj�	L�/���au��R��������7.��u�4��Xp�X  $���"]`���I�Y��V����U+��9%V\�P��,���EaM�Mp\zh6o9hM�2����~�V�N<�,�t*���o��iY�'���;AW���4f+���N�Z�"�������B.kͩDE%�ϟ_�fc��G��:k�òHHr^�Է�7�A\�u�v���GA�n䣉@��r�/KI�֑WA�"#��������ƴۗ��B�WzC���5MW�Q���^�7���{�捍b�c�+C���-QKf��=W��Ua���P���of�PB�aܪ���CS�����r�a����tA�C?��$���M��5f.'O���0po�HM4����߾�h6�zx�d6Pr��������Q��V`j�v��q��I�|��^Al��7y|��2��3����_�57*^�{���O����Q�Le�(]v���w�(�+(�{RY�D$R)Rcӟ`�zT���'�9\5 5�}�,h�B/�?R[����0�YT5K�{�α�F�D�D^з%6d$By�z���Jo�����-2�N"�����	�Dr�?'�1;�[�A%��v������O�`\Ͷ�>m�Az4+&-Z�aV����6�H�2�O�D��
��|�9�D޸}˟��&�K�>͉yź�4�`XV�B%o�"g���L����Gaۻ��%d<U�����)��c�䟼�n�UI`�h��(s_�Q�;q���E�5�fhC�:�]���8'�4���f��|��D���o��)�Ц-����=��<�x1:!1���o��O�d�;=�\��J#Yn�1�jF��-�'���Ӄ)��2t��|iX�Eq>�
�&�v{z��W�,Zo� ��!k3�T��Fhݽ��^�W �,[�n�p�&YEn�8�j��̋U�'�E���<ab�0X��M�ϡ=N�����-q(�@N�9�Xz��w����<�Q���݊���G��=�Gf������CG�������Q��$��ɂ���}0�_w�K��;K���}����Z�C(T�7���ۉ���<^l3����JPp�!�]af�x"�F�����O}gy�Fν_sՃ�k�m
�
���>���y����Rt}�؍����78�����\���͖BJ*T7�APѠ�p�f�1�fWt2�.'�ټ
�2���\�M�����]Y"�&k��#��6�bǵ4������M��x�w��]D>��f},)5_�W"�jp��"��`=�m�17�#׍S� ���BBf-"��*ϥ�ت�9��Hh*1d�6.��Ps����o����pqgU]/��ˋ�rLs���=��4�>���o�(����P6��R��܁���1�f��"r��a�ΤgBw��p8�hD�%�
�%�Ktc�a�����P�7�[Ej.u��Nb'�A���aMY��b�\x��&���C�ʎ�u�p�WSy�[z�8#u�<�t0F�U�Yn�1�n���k�k�M	e��;����D�4����`-����^��9G�EW��nI�����,�ơ=�䏚��q>�^aI�ܖn� �{�p?���E����s��z;iMoHf�~��i?��Ђ���	�X#��xj��2���)�{�S~�I�?�S�Cf�!{n(��+I�j���|�$��[ە�H�FH��y6�7.�i;#���2�`������LTv�M(��x ����BA���h��^��ީ�����o�x�+ā~d���^�\#�!�k��Ҥ�2�����}���[����"��1�WP��������)����"��lC�X�U.V����b�d? ����H�Ѻo���ֽjy�I}϶Z��%t@�7h����^���F�d���n��	����>ߞr�����T���4)��(�X&UY�qA��^���T~2��,��y�Ё����WG��0Î�qs:�-u'�j�b�z!���D>�3���k,J��^^}@|c]��p��N�gt'��0��7�̃� �,hQ�H������IVn]0���i+���{	���9A����SV�b�����Iأ�>��Eݏ�Qt��们)���\��q�"kIs�W��)ǦcU��P01#���
� ��A����`��z��5�HهG��t)q�9�hvDW�o.��� 49��!hqj�n�Qv'=d�]y����dĉ{��c�o+U$�b+����y���[)�h����\4"$;$a�3���R]�ϝ��9���� Ƭ2R�5�B�v��!�(+C�9�dI���S�죥�8N<�Uh��
n��k��p�;�����.P����y����e �TF?�skܕc7'-��%�Z�;��_�5H���5�6mC�����姀N�%/�Ӱ���X@<	0c�[߁�6�dEعJhKA�}�ɉύUgԀʅ�8�f���CE�!r_T�<����QX����
��B	R���I�`�j���z��N?�;,��̱��ξ�"3*��t(���0d5Ks�9
����C�cE�	 3b�3��������wUz��������>%7 ��q�.^���n�nv"�Q���?�%h�A��Ƣ�n����Br��H�q�H��������q���f� O@��Q�k�/�RN��SJ��ho*«��=������2;+���ʹ����<g�˶#L�Ze{�FG���w�?fƎ�CA8VW�@�D*�z�h�L�(��#O ���u�>��ȇ��BjK(i�I��$�*׭�:�&~iiWK��U�1�Y��G�
];�E�T)\��I	�(����Ӑ�%��&��:j�*޺e��Nǭ�0rh��">#��i��@]�r�'["��v�p�:	3�CH_�$a�i]~k�,����a��� ���U���N�nu���Q�x�2')�;��B���B��W�U#�_0���`ݿF���η�qQ�L�f�!��EӒ��k��`����0l4;�W����/�+�[���y�-�4�h>�F�t�3Hnn@�T��}_&zۘ�Bt6���{�I:c�8
"e3�ͩY�Gup~�)���/ȴ�T�Pr�*	�2�>��B���U�����8 �uez���x<�B�m'(�jz��|��l
{�!�1�&��j��w4��	,�e���u�H��}J/�^rZϷ��X��Ɨ�� ��@��V�e��fϴXz��]�IK�&�;��<�T����*4#e/���V�]���g:,T)��r�@(ўL2@�CQn������1r�����+���k|�ƹ�*^K��pJ���k��27�%2s�;��#����C�SߤI'�n��{�h܉�����(c�� 7p�����ffY9
��s�96VDlS�D�OZ��y0���K�-Y�ʰ�"�S�\��"���df���]<��|�����I]�Q���6�� �R����猇� nh�Ȓ\|qB��
IR=�&���)��nFQf�엢�i��3�U7����5uJ%���&tU喙�ƔP�ɡ�_�(���FTY&��џ\�mO�f�
0��f<|�}��]�,<)�{.A�S$�e�|�*�	�����
�<)+�����OE$�[��S��B.�k�Be����'aq���xݺoʎ���V���zk�Tg��I�`�:lAB��,3,'� sMj����i��!��l�=r����0M�w��5(� ,�*ӳJ�b����W��Q^�ƿ������m�Y��.ȺUI��u��$��*��{&�,Y�\����Gks蛺�s5��݇�M$< ՗E�6�d  ��hp6��6O�+s��AVb ȓ��T�)��0�ak.)|I(v#��9ΦI�f�h�����ZI6�3�'9Y��h�;_���/C�м�p(k�I��m��E?m[VS`p*�\s�ѣ���A��E��+誛���|G73��� �v,2!.4y��,]�q�%v�_Ez2��'ԉ���ĽXH�fX�+K����k��@|No��ˣY�5\�K��{z
��Z��ȥ
L�2� 6�&�f�M�|����	�t+�b�ƻ,_��C`:�徇��e՘jx�&i�а :<�A��2��X.��jkO�]Zs��4q��Q����'x��jK�֟5� 4���G6;�R��Œ�7x\�5k;	r9� �D*� ��%��~.��*�Ų�$%xM.���V�G.���)����k̔$�YlJox����u{��c)'5 �s�����>�G�Z�*zy�a�|t��-���9��$yڬ���,�@pon��w/�#_�E'�L�h0���P#�}�]�����#�d4����Y|��+� ����{]\�[R��h�ȁ�	d�	qV����m�4dI�5�Ͼ�����������ѧ�_�b��t�ߠ�~��JJ[�M��p��ޘGlV��3%����Iq�oR��Z1������K���J���1c���J��t�P:�?Q#I����bT0E%��G-ȦB�r�x2n�	"��q�����&L��UT�GR�TAc;�6�N��Bn*�^���J�R5w���9�u�p7�Ղ�`|b�([siz��[�s޸H�8���`�P�"���E6���ٙ��	�g
g�+=��QR29�Q�M�sWВ��]�,7�����G��&�-S�c�� _i	�pWi���)�XR9�����?��pPQ���[�"�,(��KH}�>�a2uU��>>E��Pj�g4�p��mr�o���M&�bl�"�P��c�Jl3hF���H�) _n�,��8�n�b��� �EQ��G|���f�S{��'J�
YͶ�r�xtL}�����<#��?�x��A��$h��BX��<����<�?=���uc���L*�-��ܢ��g��=_����P�>�>X�|�X�j��R�����s�~����©)����V����*A��C�h�j�E����w����J���R��jɔ��B��Ta~�bSS� ����ն����xT0A��b�JW��g�f�һ���%NC�whx;g-�ٵ{V�Ѹ-y�<(��U�����/�:!C�0 � �~ðON�ں�hlf���x�ֽ��9�>�+��H'
��ꝦƀU-�Z�	y�Fh}�1�c�g�� ]4`�8����"z�i"UWv���"x�M��jT�هah$��.�IW����r�#١4Խ�Y�h��f���i�|�c1��7�/��;jm'�Qq~�F�j�D��;u��T�֕X�����oĞ���IV=������:RG�P=?�]����~�I5��w�b�P��.��z�V��=�!��UI\�\����<�ǀ�z��4�3����s��d�⪣7���w��Ὕ�t�]vj�bR1���~�RB~�
��V�>��goe�|x:�4���?�����+�<p�V���'m+�7&�� %�`��-[#�ʵ�x�����ۓl�ޙH�iW�x��>ڦ6��_�(5ó�<��*�_�;�w�e��(/!�e��`/]�25��#U�*�߄�HI�;W`@�����<(G&B����� �.{[���	$���W��+�r��3�/����J���:mh���Է�)����ߎ|L�s���t7�� ��z}٣zgd�e�Gݭl�W�}0d1����m���� @%�8=�:�%J�<4}�3TԘ��z�?�Oҁ۲O�dť��-6����x�-��/N����'�U�-/h��E�z�*���p�"��:���;�\��P,?��s��>�dS^�6u��&Ldi*�f0A�`<�T��1Xx���V	�>�|7�@�M�M�i	�k�A��2!_���;�|��A0ؓ��^g��7�`��@����e愞�i��kM����[��������T2���Έ��İ�%�)�?�Ge�}�\t�|�
u���5���b�ȘyC��!:��˫L'���s�}��ҿ�ަA̐�u����0�9�SʌT���P�;y��׉	�>2�����.�0swT�-��a���4�+h=$�ࠒ��:K�js#*�c�E%���]ߞ�S��|��k*]3�E�<g"��z1����.Cy�'����]c՝�}�RK��82�,ڶO�O_EtJs��<��IOu���r�爋�t������X��>3Qݖf$�Y%�*�2��:SkJ}���`!���T<OK]����p�O}3�T{�6�>0	�H��D��4֤�!@����4
����d������)�O��Rq &Άw�>�$����3W�5!�qfc��2��V�=Y'�ٓ���_��S&��`���� o�^
���,
l��h[ٛ��B�]��o�
o�������9��N%h�<�U�����sƚ�]��(��<:k"q����� }��Ͼ'^�S�U��-5�;-��\(�ܝq��`��g�m�v+8��)�X}����/��wK˫�����G���{�t= �.EM�]k�{�����%����wnb�n���I[�̏��ePp�u�E�|.�{*�w2�s��? j�:6�A����-�9�LB}�2$o��X�!���܈P��X7��D��u�<��������J@tH79� �<-��e@�}X����M�(�`hUR?����ˤ��53?3�2l�&��E5�[�h\Dxq��3glx����0ia�L��m��C��3���QbѝZ�:O��S#��iA��~e�~�YE����`{�T�f�G�ˌ��lֳ��y������4�	�G��iGnt���wb��q?�n�5����ق��H�f�ݹ�m��$p�T��H�#��3�V�i�˧�q�� �0b�p�a�j�7:Xt�Y����O��gr.������:[��I�<C�ե	 nb���߶4	 R
��P�9S�ZL�g;f�k2�Wj*�����!��.Et�]��BF��d�����sg����|_��A�
��m�����¬)���F�Т@�����$Z��pz��g=z����A��1�T7,'�b���Z?97� #���g��!u��>�����	��8:+����w����a t6Z���=�[u6�b�0�J�Cu�!�$S�G�WK��Lb�*z���gv���qn�4X$6p� ���:�S4Y��s���ڝ�����G�I����k���������6�F�-��b�}�UA����2T�����?��b���t0�춳\�w{�5�[y4����|�����4e�&��ǹ��LPXөO�5"�I(C��n+7����-����������?���q�j���ϲ��B����~7^oà��C�Fw/[�� Qx���W���߿OFD�9��>_u�­z�x�y!�|3�Q��\'O��#��<FMt��xC�r����@�Y���5�YDv�p|����5L�E��C 7�xbrL�p�d�J���|�u��J��J�Ʉ_aH`��J���?�#/�?G!KNBx�f����9�.� �А������ۥr�h8�Nh��}��_]�7��Lƻ4bnʇ1�*�is�Z`$b���^����`�����8�~Rp B1�)D�x<���c���vxڪw���)�N�+ћZ�1�+q�{K��tg^C��݉z���L�S^��/���=��-,�m���48�6G�!Ló�c�n p�Wy%jԤ��!�u�����N,�/��h�eԿ�*��;�4���pم�Ā�-*���t�`�/�M�����_��E{u ��]'����	І����	���΄���B��<��5z�p�����C�C�Z9��
�w]\�c)�D@���Ei���+نjc�@ڮ�������(���M~.�B��J ��֓~*��lP]�s�Ŷ"2�,cr���Đ�4d�
����V�L�lXw�*�R�%n���hE�8[�JL�m�Y<.i��lZ���2���u�d�̼�>�(N�֥n�u�uW�,TR�6�9�G�XZ7Z����X~����"!�isAӈ��A�Ř"Hw��םɫ���tZ
8�	D���$Own<b�ֲ����B���$��_ :���`{];�ףx��Y��>B	Q�����A��|d���G����n�^ �����%C�zPZ�|���|�fTW�Z��@ԃG��0m#��aB/�6�kc3a!R;���RM��Z���旖 ��U6V��}+�qS�JM�ݜٵ�|+W^�E�
3M�EƷ��{�����L��ˉ&���%�'뉄� �d�4߀�'�"�I(����@��1�4on�L2!<vK[%���FW�8����������D0�.�/� �=H("â)��J(�y��)x���44��\d�~1����ȭ��(��G�]r���6h3Nq�ygVG�ׯ<����=/8�ҪFظo��D#�� ���Vgh�'��kh]�u��R�0B�j�����ؽH)!���lP1Umh���9A9��p;΀�O��o4�Q['��s�@����_�{��
tP��UfP���h�e*�#�h�r���eQ�	��-��?�%���0�~G�c��ʟ_ƴE�H�A�ٱxg\���5�r5��h���!r�N�F�{y��0F�~����'>Q���^��	��kZ��U���~&�͞��Y����x�����l�؁~p�K0Mq���dJ4TҚ:9��SH5��B�"$��3En~a�/8vt#	V��d��nl��R���Z�a[0�k��I�%�|ZmAr���!TG�V�}V"��@����p�>��j�C"��P��g�X;��Y���t�N�	ܨ	=���]�s0X���}�VNc2�y���U��ىQ�H}��OA�
l��:$����OS�ޥ�k8�>�hk�� ޝ(2�K�>�*&����?�v ����Ns��' ��h��!��ؽ��+Y���s
�r�K�N��9�I N}��y:����'�VX��Elԛp���֫�>f����U�-�)?�@>I��N�RX��ȓ�T%�q2�Z�Ʌثjko����~M1-���~��5~�;�OC_,KdϮ�5hJ���y'g�<�}�Z𳘨H�*v�zn�_fI})h�g-cw�ɖ�|�ɯ�x1��~�y:>g@�_��3��������`ʌX
�(����:�s){����}$2b��6��:q���χ���#�<S�`u���s���h,�	f}�r��c昅���b'QH�dh]��F�FU���Y���3��A\��
��g���j��n"��*-wԡ���1��������w�.ޓ���;ύn�yp�qm?M�+�h?�OG�Hm��D��re���UnHb�)%��/���w�bh`gʅ6;~y�X� �C�{����?@��kOp?ʤ��EXc���H�����{������,/�����&0wa����l����G�w<����D^K��5~��J�Y���Tr�DJ�D�vMW�?:�]�|���b��>+._��Y�筯\��T��@Wn�lH3era�;��S{�KN5^Γi��g"W�f��������I��yLBCr�z�(�^;X�QC 	gtr�o�Y�=2}�����E��Lg5/�����f����0��� ?�αf����@��p�oE�
�p��ԟ0�����ۜ�{���n���:��������U�EM�5�/uY���W�d�����'74Љ�#/���⿷�3K�涢�����^�n&��@�Ml`��s8�	��k�w���|���'%��@KC�3�Q�x��.�x��~ �W<��Q�;=�]�h;16��W�APP�2�(���k�k���������A`�K��>4a��	�+|v"v�}�i.ߵl�)���B?-+M>�
��l�VI�~�*�\�"n�iwn�Z52�����
_�����'\�x7�a��;7���c�t/ڜo����՟y	�7z<[1f������n!�LnJ=ʆ��)�m�)��ο�n�S�����fd��#!�߱�َ�D�#j5L��C��X>L^�����9
�� I�lJ���PGk �-h��	���5X����/C-����~���{ ם������&G���4C
tH�
��uE]j7̗Vl0�'��T\���<����oF��Ƕv��K�љ@Ԭ�]_�9��hz]H"��c���vQ���W1�0���5�`SBj;�$z䒗e7�stO�Z_�#��(�2\y���BGoJda렂�o���R���E�-���p� t)C�`ʷ��>u����[(��V�7��j@�őZ�ixSY$���C�:��bh�bH�NX�+��Y� ��i�\&���A��d���NW�siU�06�X�B^���xp��Vr��^��Q�G��o���vS�.ۢh��*��7�4�5���w5�����&TDe�����';i-�e����|RV�d<e�i�����%���M�L�	�Nzg82?d�#[y��1�=e~�>���P�X.�f��oH�m�K����C)�����3�΍d�j_��;��P�S���&=�����]Y�qX��1�{��Ѭ��!�Q�a���N�XX�b���Q��Gk��%��9�P������!^D����>�=
M׀[u!yM� �I�$��##�;0"�mt�2�l/T;
���ӸWK
~�K:����s�&�O#���~�Ԇ3��� �E֐+\��i��MOS�Y�z�f���\��_8ݦ�O�������%� �m�!�d&�{s�m����:o)yz�̭N��V�e������f°��`se0�5�����oT�f��ۜ��	�Ԋ�d7 pP�,�p�����A1�yź�f���h|�wJ�ڙ7m��r<5�j��?cz7�Ǌ������/Lm�����P[����5�,��bD8i�^���s"Q�L$��|��;��pm�?ʌO��0�ɛ;�b�P����@�;W;qƇ܍���3�k�>��sI׵a���W�7M���#�dX\Hƛ�2�f��b���5����i|��x�}!�*��� QNmYh��?�ϔ���q��|KSr[�S�&��c��E�Ȣ���B�~�#Q*���H�	����Ya6��I�R6%5��1U�F��m�6�+�"Gڸ�e����ɤn0�WZ�g�����;�Cz��,��I���=�|C�J�V�ʋ%_ى��a������ֱ�����\I��-"����% (��=�;��H'�|4᠘4i�'��Jv(���r���%`��4T�NMf"�MbW��6���%���v���L�7e��nB�}Ț�*�C~HX�v2Lp.����	�g�L{��^�}s7.@�z�}�#l�w^��d8�0v�Y=�i�y2�{mn����`n�L L�+6�4�+6ǐ�Q����yؙ���uuԇ<$K(�$Z4#�ٹ���R��5��U���#��0yGD�L֨W�q(�Â&��-��Y�_�2����b�@�.)B�O:����ʠlK�Q�<?��O���y�V;��b:��@���r���[�ޑR<����S.����ݎ�wQe��o�4F}�T=�99f��&���	�(��.���4���*\��{U)�쩄����;z��Q������;Zo��	1Im}	�j�b�f��C(P><(+�����%��p����_����o,�`�oD�Ү���d�+<���@�o���+I�Ae����΄T��`<�Ow��.+�)��!?ϒ�Z�ђZ��q���� ��CK� �;��|at*�MΠ��4Q��w�y�3֌��/{�e[��}�{���A��h�������/�~)�	���4�B=jZv����^�/��8��_kQ}+�Baӹ�	j��8���̧l}�3���6�e9 YJ1��v�!������\U���|�?��̥��XF�1Z �1��Օ���*דEeg��|�tm�� ��RQDʌ�E�(8>���Ssy�(8���?44�2��S��=G�%<���%z��}�p�|q�1W��u�Twt���X9�##po=�TjGl�}��<��s����r��u�KM�?j��zB�S;qQ�i�\�[8)�Zܴq��CAZ�A������~�_��eak�L�ɝF��8�/%԰��N �l��"�%�"�(�r��l�����.@������g&m�vD�,��
�Ro���0�"	&�+��âʡ��^��R��IwB��ιoc�_1��-D�E�#x�}�/�S�VUk���j�x1'Y��A���$oN*�?}�@9�e�=�0�����0�w[<\D�P;�w�	y0�{�šwn����v-z'_�����hx�'������s�[�w��] ��%��E�Iy<�
�@kɼg�\t����3	R�IP��+D|��>2���?�G�Վ�.����N.��k����a�B�8jyL$-��nW��m�����%�d�!�ڱ$ve���ц�(�XU���d�Qq�H�3K`�
�f,��Kff�ૼ�����k==��ڥ����β�NӜK
��'�(�;+l��O,--����1Vj:7�86�dB���l�kd���f.�k.����0�:��3����D`%}��/�s�����+5��'6<�n�S�wr��29�N M��iN{����J�HvR.��}v�;Vʃ��w��q�מ_Bd��4Ý}��{���`]W80�!s��#���7�x��TT�z�����D�m�t��E����mftn<�iC�����̮���}�����3bPz�&UP��&Y��Q+�bʿ[J�	?�i�L�B\k�f�D}�n�C�X�d�����,/��S�4�Q����4��W7Ux�"���\�ޔh����m����%y<�ɳ���.���JN��i����>?�ZOR�H�[
1_6T�t�(;oж��k�[r"}���T)������Y��]����@u��6th'צ�̥bgc��Ggd��;3v��zR�J� C5�,����ʪ��W�Bp��ڝ��#�@��1�U�C/43���3Y�l���Z)�G2<#��3������<|j�D����W|k�JU��d#*�S�<�yX�E���GG��sy�*��S2�<9 $WRI��7uJWn��9D�{� Z�oyK�9��w.fZ:a�MRrM��D��+j<�e�%`��2��m������҃�%H��(��Q�[���wN���&�ʔj�,P�4ℊ�**�=4�`vmd��#��q��Yx�4x.����+p$v|USUƔTt;���� ��&4u*FUV��ٝP��lxM9���?C��N��6?:�1�_�gc��DP��Ջ@im��T�[a�����vS+6��=���>��0̈R��=.A�XNO�+6$l�ͳ�˂m��i�m Nx���s9mu���М�cR_��s�iO�!�=�%F�T�ɘ�~2D&��.�.4N��3o��ǹU�4QN�D-~Ay��9&	�𧬱-�Xm����ąI�(C�r�!��Ǳ�͓�⚲�R�n��
��/R��:��[�����T�Y� ;���p�3(��e�j��� �ԍ��Or�%k�Q��[�tCIt����A!}?fƩ�7Ҿ��5�]�QY;,曷�]���'�4!?/��"��_[�g�#Kzgֿoi�NJ��	��� c+��^�?֔��+�����R3&��F�c����i�+���O��"�n���}HO�k->���b�49�4�Cf��m���F����W�����V+Rͣ	AK�`�G*�f~MWb�ǣħ�[T���N�x�������y���#��X_Il�&�u�|�e;�\mx�:�%=��XZ|�e��@×��m b.�6�?�4?��rQƷ�|�Q��n��,K=��tg��ZA���gj��Jʁ8�q\pʭ��y�z�ni�%��w��1�h�;��-�լ{�aFw��"��1xh��(���l?N�a�zä8Qy����x����k)����j7�7���{hS��������m����w�c��+��C¬��)1"��Z�(�6O��,��I�6|�+ȏ��X�J�b3�������gH����)�{>�t��Q�����p���������`�@_4��՚N[	��s#�rŎ$�}��II�F��43�"�r����[���ɵ�B��}ꇄ��J��g�Bd��SAM�){^۟�|���6�lE��}Ƒ�`�A�V�X�qB��E���OMg�+_W����ׄ=`�b�O���	.f�?��<���qݘV?�YA��4"؏����<p�8�� �.��1#��C�隐�>�������DM,z�ϗ�f�Y���l��)�@p;�à,�sU�ݺ'��;WF�Ơ���K��%�����;i���)��uc�Exl&%�oϪ/�`���_�5�k����\�bHZj�~g\t�C�I�w���w�!���R�jjj)�U2��9�rv�`�C��ͯ3Fp�#K��v��2��E����v�)�V�q�XV:���x�N�w#��I�j���X9dW{���v �	qe>��+�����%��,iwR
��D�f�Re� �a��d.����~���UQV�
A����2���/-�MP�s�3IJjtZ�-	��6��F�ɏ��7���/~��T�7��������<��R/��r�=[��:&���d�C,u��+�*Dh,����+G��d�RH�8�p�(P^�L�*P�|�6 #g��%b�`�l��R��H�M9�YM�UǚG�X��8�ope�v�$�P|:��kk�0���_y��j�O�x#w��(�o�q`.�.�;%����W��������h�e��{1�Z�.���)�����M%σ��M��c�����e��M�:_��LK!�[�����il��Zu>�	�X:ė�\3i6����
�f�~\���h�3�n� G�Ĥ�ˌ��Dw�-[�ķ2��X���%璾� �Bi��\Idt���^��{���E�2ˣ!r������>v���$B�t̖W�J��Uhp�.$��1�H��K��s�\�МZ ���.��	{ިY14�ݺ��������T/�g��Y��V���� 3�|�bG9�m4��R�s�ZPS�;� V��f8x�z�SH�Ae�/�_#j�XI�˴�H[�.�`^~���G}��ZBY>Z�r�"�j��)Y�0rG�ra
~����K}n��`�og�t��c�\zs�]��Fl���d=@Y�%*�3��h.��k�̮U���m��`��[aM6})�2���r�R���79�b���3��0՛E���|JN���㒉;�K �jg���\zQ"�����
in�@�Q��jl�*�c��N�x(9�})T�(����ޢ[!����_�+��,�0���:�"A�&�u�`��MOh�\�N�^ۿE0a� Ö?U����ǵ��@�|��"D��q�gH0�-��v�Wb�͓ђQ�Á��zIT!�%j�?S,��!�j4��0]��p���n1�ތ!��f�����|�9x-�  �r[�lD	�u��>�N矎�I�_�1�\nM���b��TA ǀ�5�z([!���p��mE�4���1	�7N��C�l����xc��t��B1G�������dV�ֺ�F�=z�|�#3U��[1���P?��Ĕ[rW����iz����Ck������6 Ŧ��#�(�R��qk��@�;R���y�o�݋@!h��X<z��� >�¯�f,,P�$j)Xg��^��'��ɖ��ީ�Ra�9~_��n8�i���F��U׏4�lJOˢ���ͼ�w��F�^�C������]o9.�{&2�����{���KS���Cx[�[�@�*����ۉeLҴ�y"�-��+��!"�0d1�������5h��	���{D�Zq�L_��|Kt>p�FUa���ny�k���gB+�Z�t�t�aɻ�3�	|ǓF�hT\Ԟi�]I�o���w�F��j�����k�%2;��?W�n��+Ԗr�	9�1�{�"�s3Lj�q:�A�a�����Aq�i�$�bL�ć�W~����/ʷ2��`_A\�0h��>Q�;����~]��0m07�5�Q�ړ���
,)�S�#��5UB�}b:�YZ(	��c|�� Ս��0�d���[11�0�����J�(�}���~���&� ��du)h�]�~�ٴa��DsPL�2���!�R���-�M�B���l��l��pN�����JJ�i6�>#.�/��8�c$t���/2ܫ��J�_�KǙr4F����$B�$������*�
��|��Y�S�	ÿߋv^���{�G�︓�~#�/�����-��m�q\(/Z��_��e���� y�u�c��9��Y��������f������3u��#ε�s9g�C�6M����\�lزB���
{�\�GN~�;���F-(��������ZA��w�̠�j�Rz�F } ���R���I�~�J��ݿ�:��f&9�B�^-���!q@+���JQƸ��D�l�h,Tk���(g�:�#e�ym��k���/��?�����ʗ��I��^�7
��F?��HZ,�|�©�#�����m��|i���P�;���Oz*I���R������!{�쿐VK2a��������n�6�]�^���&'1���ز`�ֿ}c
���z���,���[w�����(�AQ�����}RBjKR�$�F�˩'Tz�G̤�_�r�>��õ�I� �����QBuP2����]}�{ֶu����`I�Vy0'�.!����b|��."eH�����.1��((6��ZPG�����r��^��Ld'g���q2���$��ڟ�?55'h�|3���;�K֩�p�I~�B$��T[����C!z0֕�چP��1$\R�a_Ȗy[R�Y��JvI��}��DX���}8_�W�^��-�$����)Q�X����"{�~��Q�`_�<��T��8懗��04�k��(���2�f�,͔�NblH�Iǯ�\�"��ة�Rm�[�6Bш���Y>�����&�ܛ赣 ڠ��h6��+��k͒�X�|������@^b(�+��ɽ��x�tǇ�*�C{��(YI��
��+��/����-f�S��Ƈ�kc�Q�G-�B!EH)8�D�����R�Z�m{�^J�5N�
�3�Hp���>	��T}���:�I��r(0��ċ���"�J��,����������TO�p���q�I�]Ws-�ԅ��/���Z�Z��sQx��3b���FҎ�'/3�D�	4-�{�QH�]�,쉲��ΐ?���BUkAۈ)�-�R�?��y��.Tl� n�;3����6Q�>�u�9�g��ڈy(�<�������U��x��|Rti��������}f��-���,MdPP1���]��2�"�tv��t3b������r���������.pBˀ`Q�����ku�W}�d��3_#���>��b o��z��Q`+�2�|�&��b�5��HN���î�9�2zc��d3-9�{���cvu�M%�Y�
�d��u��e�$Q=��y��a2����>ڽL��n蔐��֖��s�!j�R�D^PM�%��icj��}�
��Ԍ暏A۵N{�����y$۠=��'���1����MN:D�y���T� ����Ot�Z.;�j�z���&9/fh)Һ�޸ z�܀/����h��N��d��s�7�:x�"3��A��W6�y+k*���]��̒� �-���!�XZݷ6?��kq%	�<|�
ey���Ȭ$�/��8�D�M��M��#<zf���2���~Jl��fd�m ��o�s�N��B�H�E0�T͎�H��z��_�Y����M�Y$�x���o���awinFC?�Cw-�=xӱ�����,8��u�I�{g��=�n�j�4#^+0^;r����4!"�-�0}A��C�*L� 	펨i���d�j���-��+r0���k�Ty���4A��h�����;��
���)��!i�L���96���Q�Z^rcԏ~+Rn�>fd���fnt)���3����a��)ξʹ���z�L5��>�=;;�
*6;#��C𞒩3qˠ��{���F�f�bZ�@��G�rY]�q��h���i{��;3��+Ni�HvѦp���<y�XZ�>J�ui>���kAv�0;/!H
D�<�\7|K1me��@� џU+S��B(��O,#𹢅d�U?�����AR��=�6ݦY?9��4/��.*l��E�͗ضW��o�E�`�+ܑ����c��--�^XgA�x�cѶ��h N�sή���}a�/��S�<�g���?���\�q�e����jCr�������3@��5A;i�~ H���S��HK)��8�d%��I�I$�P��s�_˩�m��0��V�����D��6^{*�%؂�*��/q<)_�:�0ѫ\�j�H[�60V*�"��n������Cʧ��r.JX\��=�kO�r.��x�#ܭ?*�)�L9������jߜ�P�N�ȂB.���b!����{3$�4�;6�q��nu��J܄��ZL?t����y�E's[������E���wHwVd��ޭbbZ�?f>�V��Z!�1��ԩ�
��d��w�#�t��p�L��-���[h��{&�[��,�������2B7�Q���!dh�;�f�l:��q�Bo�'*�%|Hc��΍�j"Tv�|K�����MǤr �ɝ��� �~�b��U�6*���FZE"A�[�����e3'>7��)��ߟOK_� b��~2���æ��չ�����i�R�S��I��`؀���z�3��-m�p'������աgV�.��L��eң�������/��N[1����I埜�b�g�]�ߺE�ro�*�՘����V��"DggZ��H̛ Pva��4�%��g�ra��6�!��i�sZ�D�,����7B���1��kݖ�
�����Z2�@��ns�Ry8~!{|�Y�{/F8�0���c��n!������4�wswn�Np^<O}z�T�(���;I�&l�;����	׶�R���<{�9�%˽���A����(�څ�^�T�� � ]�1Ʉ�y�A@������ �3'd��mL��Z�R�����±��)Pb���'�9Ճ&��1{�����&6��Kk����n>Q�3��0��؃ױ���P�:�7��F��e���z;�hP�eIҧr>��]��YXe��`�{ȇ\��fQkH��P ����X��96�,� ���X������?p�ef'�\�@Cl�[���G�1~�=�M�*eE`����e&��bϼĺӧΐ<�'��K#����. i	�v�
�Î��`;�^=M��Bs�N>y��׉]4T�~�m���H�?�rh���}�z��=ל��3Q!D���;�3�����֐0���f�Q��-��H�l�C7�W��¤�t5�F��B�ú~i"=��ƣ��\�2U��.�6�g���J��N������ፑ9x� ��o"�܄�~�4��U_��(�HSk+�`!�Tap���h��g����6of�(�z.&̷Py�2�$r��/h�m��<����2��<b����)����-oB��n��_�ޕ�X�W�lĲ#�S����p��<m�cӻ�\I ,�*�8�0��
b ��O5{R��z�����&B�j�<�)Ue�� �@"�R�I�_�^t@5�Uy�6������s��_���A���l=P
�]S���w��**��0W��Zch��B �s�� �����1��ӒJ<N����B�Ҳ�_�`$���n=F���^va�:�R�A��:��I��T&��lTV�7#?� ���(��`�\<���fW��?0v"���y����;�:��H�����{�����3˳#��h�s�ֳ[��8��S$�P�7��(���)5Z� �3��z��X~�/�X���7e���G�	ħl�$�' .O���%�)엗�}D�xt�j�'���QKKś%�����'���8'�t!��[]�Y_���X粳�ݗPݱĿ>-%��N,F�%��8b�~��yg�5ƶ���Y���tC���_���N�"����+�|�UR�Dy�~���/V_"G�fs����í���c�'F�Z�"6̷6��_]�jr�k��*~�`�ހE�h�Z�0W�F�r�_�$���K�µt�/�/�W3�Ά*���Q.@�#IA�8ݎH��~j�#���(���&Z�~]e�J3�}Hݸ�կ��m��h�����*�g�]�����
l����p�S�,QÒ���nn��'�a�e�L���|n�@�i�-���'�vnj���W��FXf�侰����<R�V��U��*��+�:���q�'����9ȄU3�v�3��)�^�40r��u��-�@�1���_dH�G5����W�W��B��D���	y���
?T3o�S]�XRV>�,Q"��"���Yz
RT�Z���++�Iv����Q��w�42Z3��AS;x��jY�s��5�q���.Ƣ��VyK�*����]����;6���|D����e�UW�19V92 UR�]%1��J&��3��.G>7]Q$���(���~����4H.�J����_�~N��oq�Sc�N�L����}>�GԽŊYˏ��+�|b�;1%�~b�^�p.B��`@`
V����-5�𕦐s�W1m�ͣЕL��1�	c�e~.H�\�aw��HH�L�;���i��-�ԨX���i��Ks�'yu���ScK����Y�q��X���j�L�%��HG��%�!(���$ 5�Ph�V�E˦b�I,�d�#:wm� L<���d<�?Fŏ�Y5�� �
�ʱ��#�30z{N�Q̫w��m�kj��L��%ګ��5sK1��&@����h� ����f
�RFZ��0x���u�C�!:Ϣje���d�w��ys�����ح��Oi@
8;Ćh�&�L�����Q>m1�d����T�)��	��Bw��]R�~6^�gu����I�x6F��&p]��r�h�cr�uj����끉)`��ÿ���g��ā��K
�<3���M�퍙-���]r��w1�R6�E���侱��1L*����I�T����_���A\���![q|�ͫ�T8r�MPN�~yy�3}ZX�xd��R��u���D����QxMO�gһ��C	�/�� �̰�����[��vӼWp��ҫO!�����*��=��٧NC�ৃ�Q���j�N��s������r������-!�_�j?��=�`�.E'\m:X:����{�c�k�5a`9�Q�/2C��������`��Y���Љ� A�S�Wkn̙��T��C��}�О��S0WzcOU�sn��n;��L�T�`T���ߔ~�Ir�%���ji��W�̖�����t&�K-�i�E��`�~9
�-�dڊ�3{
�@��'�e�qE��)ĻS*�5�UI0Nҿ��¯bD� ?��6�!�>�~�#��(��l)�%��|0?�\�y?�VF����H���9��S��r����3"��\KZ�>L�n�k���M��k���H�� ���z�x֥��V����r��O��H�-��ǵ�EG5��6�`�B��σW���9+*�����w4(���`��?��b ����,wǩRVw��nr/��[��<.�
\"3O Ņ-K������]���K�n]�*��T!B4\*؂Uo�9�(�&+F�7u���	������tȱ���������JS�"����dLU}�H�K�P���1tl�7��|�L�d�,��/uޘ��F���Q5oߥ�fS��Yx��z��@����j��^�]���-���eQ0��!"��5%�槿p��mf�s���g��洔:V�o�|��>��ᵖRi�H2�A倁��%���v:��Р��yҼ���LT���e��z?Q��X��V�����=~�`_��n�	y_��O�X%�3�fM,Z§����&Qb�����^���=�	O�Q�~<&%ټ�:1��`�u�VV��)���|'�ո)~b�'A�L��B��s]���/�%|J$�
��2�|�j_�"2e�b�p%H��DU|�*��s�]�Y�%��J�8��d�֣�����1�1��P�	���vg�&�5��_�����e���Q��%����9�� r)�J�m5��'�R�BP�Hu#��l�X�1J��C$I��Lb!�t�HO�z�>�����-)k?s�q��o�d�	�%��s�[XC��ϻV��~?�vp��u�l���Ю�y�Pl��Y"vw	�/������[F�`Eˎӄ��(�X
`4	}4�N�k�&�[�G<�@�_tX�q��~B@�"�0�gL���� �2��ö�q��u� ��u��f�1D�f5��K�x���&�W/=�� ����|�v�n՛�.+�@V#, n�X�	����xk�湏�����qj��;�=��1s� ^�p8��Y���`�C���n��1���4:�<���f�m~K������*��)q�ҩ8�A��n�eÂ�ɫ���i&�=-�Ӓ0����o�.$�����/���=G�ކ_�	��L��[M'�8/Ig4q�n\XE��}�zw#�B�C)�têܳ�zzGl� nƳVv����a�'��}�
���#�����s���P��3� d��=����A�9�`"��~8�)V6�!9�W#��e���,�ύ_��#
������K������\+ٗdO�L��	���� �g��&���Û�Ď>A���L�F�������-&to^&*cH��.)ڪ#]������#5a�=R�/`�Y7���wa0��xQW]�����2,�j2����� �8ЊO������R��p�:�>Ä
�:��%�&��
��#;!�ᒛ��&�2�S�1���}�%ӯ���M��?I$��4���N)\6��\��S�*����4���U=3��%G��:�yt(���8�YKUI 갌@�+��p"��w���F�<�lȒ�)�DW)7�AwMEK(9����x�:��~^���}G7:Lʈ���p��oG6���.8�����Uni6rKɎԗ��h������X��ba�oڱ㹝���k�tDT�힎��JrU�uO��_v���^cj'��qz@O���[L��(�������\d���/�D���¥L٪� Q0���w)P���bQܲG��蜼�	��=��t<Ǥ���0A%�J�N� J/�E� &���8�0����:��M�_�}Xp9x\�h��d7ݢ"�?���A3_�$�=t�i�Nrj瀮��T�z],�3;j ��;����N�ĕ��}�W�úi��ȋ訾��M�64�Ϸ|��U�����Mί��ە_<\7�h�Z�`��.�T��R�z���A�ܮ@a���e��&�8�ґK��!��k3����v�9�l�ֽJ�[���r���jЫK^+�[�'��[7���|#*��ͦ�+R�c�M��N�.
7�0"pr��bC��:j��۫���L��@
UЙ@̗� ҎC	j���!+��(Ȕu���!�����Y�s��t	J����LY)�A�eސ��.Ap��8��a�󨡇�`��i#�{,�F������b�j�A�*<��^7�T)���70ǡg����a(������fߑc�C�J=�+�j!�:;��<��\ �91����:w�)��M_�0��]`�[cw�G�M���&�9Qۓ����8z�i�g)l�7z:7�����~~��>��u�m��K�5B#LԊ.{������(�������8��@x&nM��ӑ1�< �E�7	��	q`�Ҍ,V��`�#b��	��7�k:BI���k���V��P=�����ݷ������������� @�\�	^��pLZ�{�@ܲ�έ�͇��/0�Iҝ�D@���>̳mR�h�� �D��(�� �R�%���6�e���s��p�e�Zo(_��1�َZ����W8Z�U�O�9����-)���N�z���)�}�yubnS+YЪ}���T��=ҬU�j�0J��ZHb����e3m�`0U��ۮ�L_L��"s_����6�xc�	�3j������ g�U疇���)�,oR���%�����~n$|��^��\����?��I�Ub1.?a��-�l�.���N~�w�n��xF&�^�����C�i�K=��>V�L�c�N\�{����9��Vr[��8	�O�G����o05�Z9�ŷ�〓��IEww!�^P��R�l��Aj�	��T�|L(��W`�*�q��r�+��c��`����wa�5 �����Jz���r���̔��"�^�uw�ĞA��Ci���]��� (���h��9��*�2lJ-����&+ۑrSM<˄vT���K�������y�
��������&T���v�����aI�k|B �RiZodY#��6]dѝ3g@�<=��X(�wl.�'V�?�FwX��Į8z�5ZuB����9��]������m�
�A{*`ҡ` �<2d%L�7?�*Vd�tU�T䌺ވ���B���/*�ru�U�v�_��c�P���%��U+��0U���@���6��8Z�*,@�`sO�A�vc�Z��jM��B6�n�q�t^Мr������8#�� hȐ�+!��1���V���Յ�0�T�W�/�7���D-��RJa�_��!e����Ndy�:ηO��0HAF�K*��&�.ICx�e�Z:d���c3頡e��Ʃ��{�;6@�'�O`�wZ-R�x������#��y�ڸ<���� �
�R~w�փ�g���f�c��37l$yԝ�~��ip��Ү��m������J�Y}��f�&�0��"��5��X�u�����UK/�h-qx�UQ5��Pp�׼����`��w�e2�6�s�&�p�е[q�@�Q�zt���kZjB�G��A����.��c�W��iԸ���B�1�j�:j������y��E=�.�ъ�R�C��왤��mh��������4�gC�5���2W��)��si9!�*>�gƴg@���\����5��J�k�r��q��U�:M|���v�w�Wޡs2�uK�؎�3�A'��@�M>��u��󑑳�i:j���$}��w�9�	�9L�Ƿǎ=x�M >��(ӌ��1�e���?�umhp�����G��l	�|�e���`���f&�-x���8eIg��3l������Q�.cĽ��3�>Vt(!����p�
�W��P��V����S�'m�W�+�5��v��Ɓ;�a�	V$
�
R�9�s�fv6��k���ͤ��3��Xꩿ�I���.
cM�t�$�R���P�/7��a�zwG�1y�!	�o���{tK:��Κ �r���_t�����X�e6�-����N̵r�;<�6���Nh�J�X��4����*��t��L�@5�t�E�iJ7=
���4���fY����܎*�bi�_q�A&o��f`|T&ϡ9z�!�ܹ�y��	�:�7=��QA����R�U
�p��N��=���I3t?�>�|�6X6�ߣ��o�̼7�5�k95It�t��+�!\A��j�m؅R��?�t�~�js��m�}�D ��=�-�x	JSJ��B.��O�mg�dन���$��K��0��Q2�>�ʡm������$t.=^j�jϔ��A9����K1=��J�@��q솺������@�S�tX5k���G��f��rn��ހx��'|Cmy��h���^V6t<A��!���IrFnz��!�+m���Tn�Df���ʙjQM�+i�l��w	�}y�g,�'9lE���� <
G:i�y��a�_�YN7kؿ 2��&�|�9���S0��cBNS��Ub����l?����3�8fiK�^EN�[�.:`� G#�t�L�C'�ft���,P��q�S�%�����I"~��2��Ұ$_�b�rB�|��?P���Z�,,����b�����|E�Qu՘R�)�w:[��1�)��Ė�"�袔T��f�<��uw9� ��#ƿ|u�9�3[X2�<(��V <���1U�tK�������B9\t+�fN�6Ƕޘ�t.ۈ�1#H�Y������?�~es����.�+�SG���ґ��oW�C�h��U��i�N fP�3;��b���F�W��	��0c���dl��6�e�論"�	��B���t�j���_�þ������W�v��8P#�2�%�[��2���ˎ?�GKgUMM����wʋ^q�}{��LN�k� y�j��_)�@�_�`Ű�V+=R�,D']-jo���EĴ��P�Wt�މ&B�I���p]Cu ��/��(З�QR�ϭ����2�1�� ����H���7�y���I�>Ѯ�8'�օ^d?f�d�(CmL��B��E!#����|W�A;�(+*<�y54��FOg[�i����: L��2]�?�-���|����RU�j��s *��q�:�	S��Y�z:��:��v|'^��mh�ȸC��e
�+ƼA#���Չ�W�MsE5��g1h(��B�q������Z)���,�=��-L�%�������������Lo3A��m�Y�I�N�uB)��!������MY��';�	��	��#��� �n��������T��[�l�ϱ�'��Y}�RsM���A��?�KY0�O\P�d�|*�+�5hty�����m5vY�봙�\�LzF�������u���cܠF��β�Hk�H
�e�B+�U�Z�;wH��T��<��I��������d
��"�y�Q��q#Qg��]�2n}�������Z��yHVJ��]S��zT�I⥁F�'����}7iyxţF!)��u������!%*�G29��@j��2�A�<T^�4�H{1�z�Ж9x�rMaT�����Qp����nQ�� +�ؒ�L=�5�p�ҫE���׋��\yj�'P�x+.�h��	�yo�Oj"�!b��6�1-`�7�*�"�|>�gMP�� �`��B_�ӽ��KW*�K�*���֢����O%V)��7��q��܇�e���V�6��<B�o��$���B������ˎ�
�g���&|�֬2y�b�wp7��J^�u�-DN�F�[R��_�0�%��|(Qƹ4|�CUKjɛ�łs?��&�c����X��u[��W��z<I�*!t>�4�^(�\_�x�T�V��;@�/��W�'�=��t���rG�YB�y�u���6�
�,
���V�h��Y05��	B�k����䪠s���B�y���?|� �"v�A�O�5WVe�]���U�m�{3�&�!o�f�#�;�:����Z���0e?S����Q!zf31�s��G#�;C�41��_-���H�U�X[Bq3����̉��݉i�rF\xE�hSV8����p���;\wk�~�<)�e܃���])��.�}�j��>9�����A�ϑꆌ��>K�]�
'>f��9�O^�(���	�� �PZv$���R���]�oz$_�&;U9�t�L��{�ٕ<��^����Q!KC~њN��8��d�1���-�8 ��+��>�84,ȑƦI��~M�wBB{R�T��8�����#�ʦ�|ގ��w�!|%��!�6b���m�/he5��>2�~�z��6U�9�,���W(Qm�p96'�V�K������@a�Ʈw�&8X35�^�k�p8r�ȍ}����x\����zM�z�t$ u�ɐA˧��I�۽�h8��[d|t�����qT���p<n/7���À�ޚ��6<Q9��V�(���,��HX�����R�a�4iד������RbLn�.��N79�r\�Lj/m܍T�\ͮ8��+p/��j��XoQ��,~�x��o�' Z�T��%.��v�َ�C&L8���q}G��"�FG�(m6��
[�����W��}O��e��x�C��͟��G#�	�m���C�JR��5_���E�vq�ȷ��P�L���'�7 z(Y�j���c3w�$@���"�Yz����4U<��Tq!6�p�s��D��:�|�t>�愃�@7�!	e]�PY�i�����B'з�k�D���t�C��M��'>#%��Я�hZ��w׀Y!��X������2\�RhCm�kP-d����Q���^�!��n�X�u���ơk���T7�$_����k0&Q����S�nIڬX���n*#O������0"|�P�2u=d�X��C5���T��'A�D��ޟ�������j�&J�-��zaH4ή�� 1���)Fg�^�c2�XX�`��)|�	��#����[T��Am�|~uև�l�C��/o��65=������B;�,G8����T:=i2G4&ktY/��w��cXRqI4#�&4�M�c��h;���.�����N��$�p�4�j��&d��C���᜿��a�����7�i�����dA����!�����/#嚱k/Ä2!��_@=����ru����4KI���(L���\c�G�9�-ʰ�k-��5�F����]�GO$��J��:ݢ�,�	�͹a��·}���� �څ��YL���K�g�v��V�&�BI�o('�"ZXY�����8����|�EN�k�19���k�6��[��e|1���*A:0�H�p��9z��!�_*��Ƥ�Mn��S��)�t�"�pא�N�ͱ���w+[8Kl��ѥ�ݱ�v}�7��������*I{��8}��*����s�Q��yXo��Z ݕvX�z��p<�� �x�t���1d&Br�S6��͎V0K�
��%f�-D��
�9�������V�>�S��	j ��_ɿx�t޻�[�՘<�
���$ͩ�m=�m
��VǤ5ۉ��8�Aē���Z���z%��	�J��S
�).G�&�����#�̻��x�e�N�UNs��[�����aზhw�n(b��^&�󷠓�Wҽ��P"ta�6v@kR�������p!���]� d���q��3��-Lk��f���2�<G�d�[\����PP
�{��"r?�����F����.�x�w^���P��@pł���b�D�8 ;cΖ�`�sD�E�+�suw듲��M��X2�Mm	����3��)˦�y	�W1f�92�eDkV�}Zc(��LmEkQ�mu+'t�P�հ;�J�3��a�����-Ȕᙦ�Z���0�T�0�j�F)�-���P���aM߂'_�c/ �W,<�=ZsDJq#���BB�����ߑ��G�J��`y?�M:-q�����^�vz�����Q��?%n�>�����$�x��-/����u���d�T�HE��Dsx~����V��V& ���d�<m��T������п��eM�DM�
�z)�ϰj�*Y��,����a��9 ��~����<�x�[m?q,��miȨK8�e������&F9�Z(9d[�{`XG�Z�w��4���1�~K~�&�/�H'h� c3�͎/��Tˈ���8E�i���d��v��862�I׷#��}Õ`��y]����4�܏�j���bI6:��%�9 �)�U������iP��32`	�Fd��	���C|��� �|
�fb1g��uw���j@����@�G�}���j�1_aR�}\����3�ܢ\���%i�o�oQ��ˋ�݆M���w��k��y�e.l�J�n}�̕ԗ����Z�	lH0�T������b����0+�2�P�������3�1��z9\�4
��S�Z��Rʘ�����$Z��P�m|"f��+�|�B�9�qX}!C�x�=/9��L��G��L6�G�j/�f�r�v+#�����"2���$9�k����tfh�kY~|��T���~R#�T�,䶛+Gb?�"w���)�!�#��o��1�E��@�	����*��b��֠��'�{��ɾ�#���h�L�IA�EY1��R_x|�����}�����^W� �Nk^�!UE8��e ��G�in^�&%[h��J�}4Kި>�J<�驉@�πn:ߘ��4�Ћ��o͍r�l����}�9P�L�*�k�g�W� Үb�NG�K�l���5�!�#��ۍ�s�����ZZ�/˗��e}E��c�g��vdzZ��B�;h�8ԕR8Ɇ��p~�f�ǹ��P�dS4�.�uV�Yy���#H��K[th���
�9�vrvE���u;O�G�oh����~�O�#5�tq�,��d������a#����]7�.�Co_wJS�n�W�oP��s��it��z4�I���-mbX�����������b�
�i���
�NP��æ�I����`�(j����C@ά�>�����rgOi�9����貕[���=�v����_"ÅY2���.��� ����W!f�ɇ�?T��Ih�5�̙+���h�������4̭9���Q�ߏ,�JTN��*aE�<���`���Y�G��6���q�#��������������殇({P�فrr�����`��>�ٿ�e_�Dk3����HP��$�L�n�j;�����<��C7�A}���;��@(�����VW�F�V�H�=�G��T�jN4Ds��a�5}�i�s ��{�f��z�t'���~�4n���A8w�g%�� ȒhD����Jp�GO�lj�Bq�v���ʡ�*�O�7�R�9�WS�B����{�>,�E���"�)���f�����H:�����9?�63
űg!�U4��8�G4��u�gń���4��#������Ω.��:ss��D�Ǉ���q�>����ˈ-��7�.�K��3%�a�h���LY�[�Zwo<�s����ZXR#� MiA��RL���9��.�+���z"�V�j�@D���X8��|ʝm� �V�W�)�{P͌ 6u�%y���0欎N,���rRE�T~���3�F�ϋʯ����O��7b^�;�g�o�� ���ׅãok[p�X��ث��jLv*3�`-��5��W;�"�@4���4/��^�����������ь��e�ye�''ow[�x���y�r@����jM��ƿ���/^�:�z
&��;�~X��Ahy2]�e�
�@-��GLtV��E���o�*J�����1��خ�p=�1����pv�WXC�0ֽ���Z��c�:���U*A��IL)��Eڋ1p�>S��0Ӊ�t��|����}�����uQ�u���"r������}4{�.��q���e�/Ҩ+����Wv���'����@��d�e�C?����D\����|t��5��mB�� <_bUq�*V��T�=V��ڌ�K���u�D_x�5q��SSH��Q��޻����Č{Y��hx)R�E��s�{�"�C�����u04����>½�`!w��)��ؙ���3��P3��Ӣ�������p�r�?im����
D����.��5β��,)R�bL�0>��22fb%��د�M��I�\���ӏ� t^�x6�͊��˻9GZ�]V\N�.�"+��VX�e��2z# �u�¾z��zb���m�tQF�E��8���jU��=Y��"a�����Az��9m��e[��.%oM�e=�s%�Z2h�K�#��[\;�Y}�	����D��a`p����S�ݭ�	y�2[7��rϝ�N�^@��vT�������]�M��&�g1������U�(|E�Y3�"�D8aJ8�Ly�*A���~��s[ �$��,� /�RS�߰�P�]�]"�A&r�� '-S��!��=�� �.a�~���;IK�����d���.Mf2��y�aZ=}u>/��-�����P��J�g۠5	��!u�~"�,}�>&�D�+b�	`7&��"�底^S�@�����Z����0⡕J����Y�d���r!��Np)a\��3I.~�RmNg��Y����4=9c271��m�uڂ ����F�10�P.�!����_�7���?d`y�oc`-��s����T�I>�(�vwYfM�M׍���Ea��"�����1�2mٓ�.]ZQ�
ٝ���|�NQ����*:j�/,�u_�h:�Fj���QI"��#P��nɴrD��j�L"�J2�V:G�D�;�[�W���ܛk���I?�|r�4��2p��2;�^$*���~�u���i�)c�N�6��D��Q�C�\��l�g��ڷA��a�u��FMoM>��s�W�YT!����ߠ�a��2�=�"!f�1�Je�ѱ��V:�.8Bg��pZ�52�}>�֛��0���m>q�O�����ټ`vX�gU�E��fu�ug1"�#Цd��k�p���ʅ+�7ǁ��b�b�Fl���%M2o_&�-:+�
;$B�6�an�V��Ǥ��@5��6n#�+4�æ_[E��Iz�� ��z���.��֡|�0��������� }u{d*��~y���&�Ng�]&��GQ>�ɍ�"hȍ��&Y_�0 �z���o�\�~?�TP�'�WB��h+��*:��KX��5�p��Z!��t`:g�=�{��3^86�!D�d�S�up)ݟ6�7��_Sx��O��
馠m ���)�`|��EwH�|���?�i���(.v�<�LX�Ҡ~�G���A
,!t�Rq�8�U�yn��I�E�w�����#�襁U{���xb���9j�t��'`��t^��?4+��,s�m��f\��GT;k<Ԃ�����T�KVep�i��Q}V�=l�-(y+_j�����v�`ߟҰ�!;��8R9�����l(E�kퟡ՘?���F���E}��ʎ�a�����|:���M�զѦ09d�=�"�a�f�]�v����(z[3�o����=�]�k%��u�8�Fe��ȐHSʞq2�s�%M��|2���t�}{7ۉwj?:��W|��S���-����j����n���Ii+���Z��a�N[�gzI���r�z�b���9q���H؆\�m�aT&iUΥG�tLwV�������ٴ�_-V�<�)I�ڹ�1�����z�a���h2�;��cc7��qp��+7
	,��A84�Q7"�����{T���;@���(<Ԝ��w�ܞ�n���e�룥'��:�>i=5F�KO��kG�#��Z�|Y='�L�`�|܁�e���ӑ+�	��R{�ň`<���Ӝ�M�:4U�=��7�S0Ri�Ԁ�gm���+/1cr�����%M!n6�Cα<8����24��t$�5�5�v�8ṧ��؜9����eĴ���թ#��(�sV��Y.e�#xbܳT�(`tV$$��p��KV�ӻ?ː_��� ��w�({Ghv�Py�FeO8+#'ܵ���|��,Ph�6�j����y5����������c. Cu<��-/G����/�uN�����o���&ck1��,���x���«�ܠ�Pn��_����?̿jp���.#���Q�tԉu�E��%^ʜ� D$���I[�q����)T��z����C)x2!ȥn�bm�v�I�;�:�T����8)턒9���w ��N���h	�����^�� M���x��ʬ�\��~��"��Z(xu�u=9��l�H�OW��%`��4v�a�"�MziŘf�=zH�Q�`�ϑ����r���1Z�&�W��ƕ��"�ɩ���H��{�������ԟ� [��w	E�Ǩq��L�~��e~͂���q��������<ꠅ�����E$��=��k=��nCx�,#�;�m�����#���,��1�8릏V����]�i�u��ؿr��܎e���Y|z,�%���@R�M�I~,�1.��`�z47z�5����+��u��oc���Z�z��.,r���h�E˚:�h�	R�Ğp����r���fv������w��U�	K� ib��a�ퟔ2�7%���iRןݍ5 A���=d��e����D�+��c���e���p!�4ѷ"U��Bv�;J����=s �{����X#q製Hk�YW&�	ᤙ;����)�{�g�a��n�/c���U9^��Շb�2T������ϊ��K�K�BK�8;ze�����ä�%ϯ���3���g���;%�=�ʯw�l[�ب��S3h��͜���\CT@N�N'�`�	p����4���v��]�4����y�>1������l���ʂu��<��X�ib�$��y��`V����f����@(�	n��X���&a�����y��@C�%��	�U�aQB�����k�N�����o��-^*���r�퓳�S8����Q�P�H-`5ވq�_(1;�+e��\���R���&�?�5d�j��H�(�rW�V�VuŘ��6z�}�*�y�Ő>�pb�a^P�2WO���Ԟ <��۸�G�ε��x0��-$�'��[�m��#��'��
��k�*�=ϧY����u��E��Ҽ]�aSp�D�b���_�\̸Ӎ�|��,�ģG\��Ȼ���)+���_�cV9[�)DK��"����`���Q�vT��c�\�Am����@3�e<j"ĭ�V��f.�9� �h����}�0�_�B���0��&P�����Ch!��k��vO5�q)ڐD�A���l�{�Z<\�R5�= �z	O�TK�'86��	��i��l��\iR��*������]w�.�o��`=L�c�c��Ē�җ��+�9�W �9�,��{jb��<ƴ�)_���Ť�b�S݅��(�l�I�4ԕ�+!-,��2����]u��	Ķ�!u(�LZ�F���De��+b�|fO���}m����l4���"%��oΧ�uܨ!t2����K5�$� ,%O$���k�Z��U&J���	�g��Z����qr�R��A�C��PG�Iu�P�q^?���@]�7����F�� A=^�FFy�:���4q�R1N&9ǝM�,A�lK��F�p?R�����R��Q}�7�-�~���U�(��oa9^#i4���H6�l�/BA�˘��=H�(�7vFD�� )*�Pd$
��z�D�5��x�_���}��U���ԝJ����(d-�)T�g��m3v�S���7�Wأs��}�3�M��Z�6c�]r��%��ͫe�>��	b2�H͕�Ǣ�><r1�h{F�"��Ft�j&R)&$��l#��RaR6����OY;�*&���+�*��`�>��;0�.�/�������&贊����Z�u#�)�y!]J�|��6[��U��O���1�Oz���+�����ͧΣ#�z�K{m�R�u[/-���o�7�4d��ʬamc�� �ºU�	̜"d�mp�Q��ȗp1U!?��8C�����{�VV�<��{31L!]�ku �fc3��U��"�������(*·�U�"�c����d���\8-��Jmf�3�&|^�k������(|�ѺY�<hI%T؊h7����%Π喴Er��zXX��8���m
�gd5��Ҽ����|Q�ȭ�e���,�>qi,,������O�B:2�?���X���݆�f��b�\_�F�zp��̺�k�N�J�8K�@��d�C����G���	[66�v����`RtU��.T咫�XC"ZU�xEq�$��b��1�LO�U��uL��gw�,�D�Ff4����@�����LG6��/��3��&�%��M�1���Ʒ�he�]LQo��bR�����/�b�v��D\F�>A��n�pY��X��(��q�{�[�!C��/����|���Crnk����n�k���]���Á@M�lu��C(���s0rXj��YR0M�����9y�K�#e���\���`ʯF'蚫�k���#�fB�_�W��䨝�5d�;fڄ!��L�׫QO�y�����׊�D���&����~����b17pa�Aw1P2�m�}��nsj-܈X�k��VC�C�� ��M�qi�%��Ȥ���94�f$��o�[���63�:J�H���I��~�v��A%?���8[��N�!O����Q���ۜ@�G�Ps����9�?c.H�?V�>�%VC��������{�!h��� ��]����t&W�,��g���U��=W�����>I�bo�P���a����E*�Lu1�"{FH/fز��Ƞ��@�5S1�����ϔ���.[cH�����=��<�3�Ң$\��}��]����	ȗ����t�y�-���8�<_ �I.F�;S\#��Ly���C_Q�Z�����:9�2�W��&��~��a�"۳��%h
��.���m��J�-ή/�Ͱ�
����x����:)--6�D{��`�#t�c~�~����T#�K��t����> �;��"���F�1d[�)=��稁�MIfV���sH�G���v2=��5`�Zt룐˵ճ��O�|`��-/��b���Y�PN;(���~0y4��xV�|5�5!4��f��{�D	�jKT�@��]7�la2����Ә��]&��y5��~Ȃ�xK���4\���!�:i"��F�R8*�զZ�Xs#`M�}p?Ͱ���Hjk�n���^�4|0���.L�
ɟpl�����*����&A*XE[�z�L��3�~HJqd�į\��:}U��)�u-�n�����@,{
�@���ah�c��P@گLn�2~g�nMQ��!�;uM%HB���� -�G�Y~���m�և�-����|]s��!�����L���\KtK�y��^ݼ�Ƞ�ٸّ�$�i�̫�6;�$
�����I�����W|%J�����Z{����PLXU(�7�~�"�sMT$���������PC*f�[9����3��e�3hr�rz��gsf���bj�4A�Aw`K�Mù��E���bEu����43_�Ř��0��jX��K�&��e�/�NW������ʹo��s���v��fupX�,�A8�6Tk�z�l>��R��P�Z Q8��@9��h5���T�8G��T����̵����%�kp_��.�9��]#V�R�	*r��^���]zf>��3 �tC1;�k>�����L��\��(`���q���ؔQ�f�^z����S�YaE�avr'�Թ�%�Bs��B�a�|5����X?��ن������2�Z��s�O���z���>�^o�k{%�C�|���<�SF���S@8���`����|=k,M"�Aژh2�b��K�nhfTo�hcv�������&�� ��=Ō�U�q��ݴQ�,����XT��x�^G��T�u��\�`~�}{1�(��3z��;��y*-g��7�蓴-.`��}L��D<9�+�^��i-�M8H��^7��Bf�as
z1�Hm`n9��&�!Ak�\	)n�UF���������ڻ��Ӄ�O�dwx��nc��LǩR/��%��-HpY�ԭ`2q�	;ED���{p�xD2��%g�{v���uY�6��#؆�s���Z�����.԰��L/k���J��`eO�؎�M)���9w���<"&W���z������3�'�f��aa�LXrFR��4��KV!F���n/=q�q��J��ZR���F^�O<��1<G��p����7S�,6 ��ժs�u���:���D��Uӵj]0��Up�<?�o������;�x�p
?����Jɀ�9_%�R�.���8�^�jxX��yB��C�F͕'x�w4IN��i2x��,qy�\�YX� Ƕ";���[h@��U$��.4�ϲ_g�^��A@=K�r"B�/Y����UJz�@
Z�۶7�+6F�P%��k�\���,3�^d~Y��j���(�8���sw�����&�C���. �Q���=��f�}�t�8ϯ�W�\�Ϗ�Vl�A�=�$~}1Z�n5Z_y��{y�m��F��Z�F�`�0������e�8W�>��D�\+��x�f���4��o�Ϭ��)�Ǟ l-�\1��1���|_���z ��L�"zG�-Vj��Q)=�(<�4�������ۅ��e�m��ku������0 �/��늋:E�7:���/~.�������6`[��r�o�+t�䣻@����]�^���$GW���3� q>�G�f��RE�*J�B-���i����Y�fe��eQ��L�vc@F��F�${�־5�X����dpF��QYa���4��G�*c�ABg���/몊m*�3�4M:�yj�-�:q��`=�C1��X�b��ƣ"H�pJ��@`��WZ]�0�3�)��s6���X��ZDqzx�rB6f�/�4z��ш]��)���ɯ�Z�,r�W��$M�,N��GϜ	�٭F
!/L􏧞�E2p��ʺ�o�Y����{{:��ܖ�\<򖎭�|�a�d��	�ѣSp6?ά���8�'J0��1��5�A��}�2'��Q��SE�SqF���'Ⱥ�Ő̶蓫>BK-�����1�aTsJ�'ۏЂb�|�z}!'!1��V��pJ������#)[��5 R�:������O����ÖytWg�3y{������@�b�µbcޫ��3]�z�%u��%J�����n���iI���@�S�v���������<2����S���K!ͩ�HGN�t��w��e��/���(5
��:i[͡����]<��f�@(_���$�(Ҁ\q]���y��B��f�حػ�w���j�s�{-��k��eW���ҕ�,"����Nk��j��sK�L��Fi#�Έ�~@e̦Vq���(L�ݶaZ6WGϺ�tHw���!�Ϋ8����ңHc^9m(�`Jb�(���yأ����ry�#���	��Cg��I���;e�̽A�R)��`���%h��7�����{T��
K�<���&�2 �H��.�Ҷ�#��iq�˲��5fH�r��Q�"I�:O��cɑ� ��pgҘ+������#�o����?�3ab�-������h����@���`�3I��$݀U�*.;�m�ϥ��K�Ҝq|مzR��b�~i��&H��x"Ϸ�e�ˁ�ٰ���i��O�����.�a�7�(|�����T�2_]sIv�i�1R��nҊ\~N~	��4���:�����W��$�q���kw�BfU%�d|6��9��z+��l�Έ>M���] �y&K����#8�P#?=��G)W��0�+��7.�3dRd�V��(f9]A�-�=C ±��;���A��{�J?F��Kz���$��q�����
p@'�Z|��#�j��1�����ej��҆�)�6196�@+�a��Ds���P���q"�m�L"P�?�J�������]t��zMS~�<m�,0G�	��ebM@q�ae���RE֝��2����S�d�	Է�	|,O��$3U$z:C�n�4=�X'[���@�i-�/�_���gs@튄��J�^>HZ#p&�P��(�����f���
9#�s(���w��4��Y��c}UA�v��VK=bI��~`�CQ<E͊*}�Ee���rNDo@C�#��q҅��j��}+iSGsc�ak�;
���e�3SQ����iiǤ(0&?�/��i?ԺrB�5�}fokdF������N���)8���I���v5�n�GN*il\�	(#�%ˊ�r��m���v���E�}��6St�06k��=�J���6��+�� �_�1��¿� \\X�������8_�&�zt:.��ny��|?�͋��h{�(3D��N��'���U���C}hbdl6�vF����eFgIw�Y�\�}h���4m����q��K�o�!���B��C}�K�ԩC+`�9@7�P8+(�(DEM���&E�	{tU�R�1�o�LU{p��)b���=�����1]��q8T��~?���8۶�k�����X>r���c����w��U����!���BY{��HM�gD��n})աA���;�����x�{���nm���Q7�k�X-�I���L?�\�_�U	�o�yt��
&�����$7v� R�5-����.�
�cF�xV" 9��&[�d�h��G�?�@[�����j�I>2�gF�wT�wWaT�?:���y֙v@��r�$+t	rǫfM��>�s\��n��p�W�(~mo�2���A������>�@#'��j�i�Ǥ�C��~�n�f�w1�]b�Q�YǓ�Ȣ ���R�=/-�Nմ�T���_��q����)%j�œ�6!����:�MY)�3f���6*5�����Z{��@�:	�Y�wa��J���ML;P��Ւ� ������`"� ���ٳm`��8��9K�\�����թ�G�hӡZN�ND�C�bU(Z{k��S"�׳=u�
�vm�?SA�N���c�l�$��#`n��+ػ��dk�}������ǷM�i��t@Q�����.�����+�n�6�o.�0��N(�.8fJ��xm(CTi��L�|���{dV��Q9�n�I��>��o��9�T��M�&~(�H󒏳R�����*"-��v5�I��1���z�Y'�z������բa�G�*��b5�[2[��{-;ۭ�7H.++���T�4V��o=Θ�5ܔE���IB�T��;�����+p3�$��> 5�"מa���y� #�p�[��-9�,/��(��-.g�,ڊf�G:�5:ami,}A��,�l.����7�p��&�5iJ߆��������N5�YW�+ٴ
u�V.�j�G�L@0<�X߰:� /7�Ό�#C��Ԭ����'��9X��"$Q@�``=��	��sG��܅eFg}���z�o-Ql��8��C�A���ڎ�������:&����	�����I�C�7=E١�5�ݣ�F��g���9b����@u?������Xl7t�����4rU�o�f��z�(�C��M��D�V35mu��菉�F�(�Xg�L^�
x�Տ�^�V����NX��	�Oi.�i�gp	B����.dM�6����1�<�����D2*�M*��֕'�t&4
�����O{~�fB���`@��� !\��:|�<ڂΖ|����?�L��e�%c-�	(����e׸Z�2��?����h���������Y2�i.خp�1�K����dp'2�ݽ��;m*�렉���L�҇?�K�8���&�,�"��%Z���(�'
�$��a/T���޷HCo}V;����e-�˟j ��.Ɠ���}M_��B�MR�>���W�;�a�d'��!?�`�N�E �M8��7���,��~�qh���=��~0Id��_*�h�(��y�I�b��H�������FLތ��Zn�
(/�}ij�����e	=���g�f�L��f�pɪ�Ҁ��T�]�z'�)�|B��C=1��vx]�ZZ��"x�3���$M�Z��R&R�7��z������n�!Y�BY��E�,jWS�(��;`��Kе��L^O����-^.�)~���A�G�S�F���;b�_�C���,� =�����kBQ�������������4��I��V�g���Ӹ��Ca�Cl���7�^!t"_[s~� W�.����Wi�`k��������!޻�w2r�I#��E�P`Q'�r u֦Q��&m,�Q����m�|l]J���e��C�Jޱ(O<8�/���K�G�gl.
����g��P{	5��k������)���Rj[�Ha�pt<\k�N����mf�ty�_<�"HFb��xc��A^�55[z6U��,���eO��8��mu���N�53U͕Y���˴���B�����M3�����T0h�I8^�"ҋ�{MG�� ��¬}����H�1��.�|����4>g;r�}�V��<�݌*/*�d>G�J�c�eȞ`�{��a��*�o�R����P��NE��f�̏�@}�z�p�����Kg����?�o�T�7\�Rjl}�Zb��w�'�`�e/�L4�v���& �9!� Y�aO�
�R�&��l����C�f�#�H�B��KR�95��gg^koG����9{������ٳO*��Xz�(m��3�C<NM���MVp��Lt�����M��eVc��m�\�E?���n�+Y{c�3ʃf������+��������	�P�_%S%�,e(��@Ґ� ��}(����-~ۡg�5]��p��oc���0��\K��Z!BĀ��խ�Z�u���	�"гVN�kG3A��O+���B.�B�a�a~�"���#�F��������Ds<WA�*Cy��'Z�'�^�8����{ �4 ���\tjY2k�w�Wm��z�RиV3�17vxc|�JP�!�u�w|2�0�_�En܆\<��5�s�����+���`��E���<m���>�쩯�~"B�C��
y�k^y)��W���*��Z\�q���B�i�	%�VdGv�9S��w��t ���و���á��^X�㑦��0��}|��\��<S��[��W�?#����Y��Gy�[����^I(��F�vnu,�}��2�`�ڈ�#,�a�Lq�RN��ʵ*�ͯ��ӏeQ�p�T�++�I�Ƽ=�*�1���c$_��{��s���_ɧ�_N�ٮ�ե����֜�kf���v�\��0�7��j'q�#�v��rt��2:�7>'��s�T�4���k8�
q�>�EU�����)��T95��Xi��@C��!�=4�r�|�ͥR�%#Ԫ}f�"4+z���p�$�<�tv~j*�g�p�1v%D
e(0�XX�l��d�ط�9�&A���a�5�1�h���o��lk��jRO"��s'
J� �����}�YD�� ��F����j����
����}z���+5d�,�3�NB����4�N*�9Ħ	�Cr�[�%8�~Z���^�`�L�V޽�o�2ʡ�E?9��<��0H�Қo?\��Q2Z�x�"���[�	�z=+&,`�D����h��`�ו���p%P$�yq7X9R2�BJS�g�<��0����t��ere>�tb4��1lY������H{���Q��+L����6�W� ���Yf7��ZX��J�Q�RmJ��X��zG���Q�D�K0G5w�a]]�&�'6+uP������;?ٲL��Й��B<�Fh��w_L� h!`�������h�\� ���T���~�"8'��Q��<�T�A9v�q*�%⿗��M2��H?B��8e�N}P;�@lT/ڮ�1�i��Fa&&��\)�+�*Ђ⹧=�'�]��K[J�z�#2���� �e���|wV��L]_�I�hԝV�j�T3�)h G��{�o�����׽�':��QS)�S��\�L�-G�,|ɗ�E��S���9���]�'	(�D6Jp�����R�;;ڊ�iޜ{�z��:�B��ใB�	��G���� n�(�!�'T��x�������C��DY���$����;b2��Hlt*#�ؠ��&�ܗ���e���|����mw
U�@�5��
fZ�3"#���V7�׻�CRU����/��The�Ѿ��O����BȟiN�7���������S�;G�S���������\2�`>��5�����q����X���(���Qfl0o\Vh��v���?|�Ld�iZtu{��M������f~dNɻ��h?,�`s@��E�@X ��D�n�UνUoSqWs%�����U�xA�R�Iz�X���G�tGKL� ����A�c�j?F����EP��������>#t�L`���iD������q\�)W�լz�˚i"��ql�W�����W�%��W%te�bwY��Yl�3#���^�NF@���j܋���sx�1KF+s?�0�,G1������6����ʏo�B3��"=-�BkKv��3eq�Y|jJ���JI�,�O-��4��cf����,�u'^�]g�,�(��ya�{�PF-=���mgb�s��B(H()I��o�LI!�m/�Rޱ�)�,��"&|y��M8o8����r_����6�]�ܴ� [d��8�0�v�3��anV��
��
Go)�"�l��+�K�aS?}՟��p���L~�K�9D��y~O���c����H�, A{+��k՟��7婓�XaYY�+#I�ʩ�-����ʷu�+�i��+|W��օ���[�
x[1�/^�	C��TgJOv�Q
x�|��鮇n{��c8eXF/�]���t�+~��R�* <���33�^?'�&1�J������ �VaW-��V��HDZS�6~s�|$T�mZ��d�S{��ţnlȼJ��%��uOG�w�s޺v�+�+��\���:��Yy�<�U�D|�o���讱>X�>#i��\�zz�אjE�Ӈ�	�u*
>��ᛂ����=��!�OtV5�����s���
Z�y�3|mB�?������7�8�ganM�)oԿ�a��i��n1(j��xk��H ��r���e(��#� �<������ii�1%:&��E"X�Pk9�){ֳ���
�#��=��\iV�f/�������Z��-jƱk�1{������)P�Yq��K��d<Vh�Ѹ����P(g���	��u��T�+���t��l�s�6:S��Q#�s�Ϩ���H�"��GB��qIOۘ(�+!d)"�[c�B����j`���yY�Rº䡅�[��Ni�6��v5s� ��8���uz��z�PZ�s�?=[��}�:��)�f�v&,Nhǌ�'��LקOUXXUq�����fW)����]$��c�Vp��q�#��cLť����#�JO�
��X��BhT=���� I���C�[��t!̾O��� D4����H�a��S�hicT�0�8��\ uF���8$~1���lY�X8�.�,�Z9(>㿱t� b	���;򫱢����|:y�Y,`z��;t���l��	���GNM�!>b�Yd���)*�j�S朤h�X��=8h���O;s�f��<}y?�
VȖ[�y(��{�Zu_�܃̡�$7�-b?8��?��Y��I z�:�����"]�Ql�ĘG߂��(�g��oq/�O9N��l�u[�3?Fx~=p�Ÿ�=o�^���U�r#'
��Ѻ
�4��zXû�_m�K��T�c��-���2�oL��	��|e&:�����g����>ӷ+�Z�/^1���m��Vΰdp,/�2�s&;��4�egA�M��pɮ�I`ϙ)���)���Pɾk��
xh��,�/6�0��d��I�����& �/×�.�e�j���>wS������Hs�ƾݢ��m-D4P����g�J'Κ��wĮ���<�>�x�8b�!��z�Sذ )6�}Xl�v�/(��,����s��}-��!�'L�B��OMP��o��},-��?��+���İ����̗F�3�+8!���/fH����U��*+���3d-\��@�R�Ed9��Ò ,�\ �y��D�;�?7"�P�x�ڮ��aC�ypp�M�	&�'�vz"�j<�]pJ���H�y@��T=YK�Pg^ٝ�2��m/{�������N��9�u�E�A�V�CW�q����q��6���)S�E��VwJ$D����<�|�RӾG?"��L6UjI���{���|������L,��:G����I�FBY�ț	�Tߡt�O�i���OȆ)���<C�vQ���Ed���2L��:��?�K�g�ڱ�lC̓<�D�s���S�A���p�ܲPJ�'
�$�)�(�6�ڨI^/���h�p,8O1z�әsy,�9%j�t����A.v��-��a��::E��Z�x���Z=���P�I[~�'�v�Ǫ�8M��U� ��|5eշ�V�lN����lgś}�v�k�O}w�?�8��wkI���p**J*~�?Fh������x�ONć�zam�H�����"A�H�{Q�3r����0���Y��t\S�u�#��r�����.��Rץ>06N(f�V�}݈� �.�작e4�y�N�O�
�Jr"B��įu�v���9�'	t�lD-�4�,��$���{��G	Z��Y� �GL��Vs�e��p0�����\�q��
b_�J�<v�����k�nL�a��QqQ����I��s�3�#�ٙ�R�^��V�3#Y�3�5��{��r��]C�`���p3�0��GE�����$QM�a�r�"\)��8�9���H�	��h�z�~N�&2��0���H��+ۿ'�����":X�R�R�9�׹�~ +���y�bDR|gVz;)�
f���X9n#>;�+�o�t
�Mr�:oR�2�A�����\u��L_(7���_!���b2�ݯ��g��8zF����������IhL��x����g)~��z3޸�������b�9�(��.F�*#�V��wB���c�̍�:�'��汆@V�؏+;�,�N2��������?�����c�7[WC�a ��>�[L��]����0�;ms�𾌀<{�K���m<|��D�J:� ��G�ro�'��^A*�x����khp��Y��ԡ;	"��	���Ab~��H�ۇ�m_?�,��Uf�-�iȈ�צ�Z�m��B�s�^v����_XÃ��i�]�
��H��'HH��#�m� =�DH��~�WQ�C�.u�l��Ⱥ�I���=��K"�;�9���階�D{���;hѤ⬵+GЭGQ�5ͧM�@HKV��j�?��\x�1= ��_�y��g�0��g)����M(����Fg�}:yR�w���n:Y�,ڲ�5 �&��AF]�־Ivx,�8;�N?4��S��0أ/��7_
#��/;���f�|���+X���w��U!�C[?6'�=:z	&3�9.z��蓅g���(s�
ã"7�d@�
����ڠg�P&E�C8��y"L���Ov:r�Lmx�d��*? �o�E>6}����ӌ��uD	 ~f�&L��`��KD�2�Q��r����3]K����|��`�!��1�4栧�њ��8�<�<����/1�7r��c�{������ni���ak�/�r÷�����w_�C���=����jYq7�����6���ch[�?\�G P��tN�tt<jM��Z�C�ȺC�!pB�`D}Я��R0ۢHIj����h�W���H���Ž��~1�̵�%���K>4���Z�b����p��{�s�%&o[d�����s�o��u��G���A/"}b,NǿXE\^���ׁ"��f����:�gP�W�`3ӌ9*��j���H񚨝~w�6}@�"��6q��r��tG�D�)<h�vWd
@��)(���:d
����d����۶g���Yԋ�}���"d&!,DP��ɭ4��Z��E6j tn��b�S�c�|!����ˮ�Y�B�T9C�/+Mڧ��l�ё�t��8��fP���@\U�P�ĉ��J�?(MXv��,t�ﲀ��h�B����e-}C'$C�d]W9�%�i��l�PA�B�6��9FaTj���+��r�a�n�@%�&BQ)'��9y<���RZ]q۪�W�k�|ۄ̐�G,�Q<e�z�E��2�a��C\=��0
��������E���9����-�(6��O]"l� c8u��ܨ���}y!�� �M��h��O�n��qݴ<�R�ӂ�`{�<�#-����p�zq�e�:�0���UJ��=6/�c��넊^FI�gԹ��:�j�wdI��&��s�R���!��כL�r.|���U�I�X,�oH���M��ͻ"n
9�D0V�}90���Y�x�XG����c��
B~b��t3RK$�E:��+�YE&�b_�`j�6�6�U���]8�?�~Z|j�L���#<枢�)��$#FFet'֯��_��������Y`���5���8��� o�^�6U N��h��)���AX�Z'���[�дIl���s����$�ĭ=hNV�(̧ʬ�9���*y߿��{�42�D���T-(��aq%���ةO���l���i�������7���+�Ϙjnw��֓Ry�˯��96ԭX;eI���$�?�;�Y1M�rd��[���R�x�R��-G/iV������1��1⟌ed�s���4��p8q����3�$�i�%�IFX�Yg;
3I�=�}_:�)�(Ը�2RU�>���3��is�H�/��m�}�-��W�r�w�p�?ߤ�QR���o��A�h/+�����j�M-I�\TGj;�N:?�u���El	���l����2��#Ѫf���w�'�<���)fIL��E�g��ME�b����`����{�A�xO�??q��I��i-��:��D&�1'z���������ő>�AK�?-�Ok���M�-is1]�Blᣎ"�V�b�_���mٳݐ#s%��"�M�n��&�U^r޸��%;$����C�ը^l����N�y��%%�u��[��k�6�@��3�{�t�+?|�aD�&ڂ#�l��m���:���ڻ+gI�$��2\UUWú�5v$����M�y���~8���W�.��Y���u;;יo����Fa�q?��-~�{=�E�{H����g
j����\˦�g���e&�t�~ �&�ډL�BYX�qmA�N�]U�3��������ZP�z��+�&��q�!���W�°6�^H�CpN���%��>��$����ɴ�I*�U&X��Tbצ��=Dv��0Р�d/��]�E�E�6�����I�hه�"��yyn�(3D���sa�ׅ�8����.㣊��x���9-���(1	�Gl �����
l1����$!����6��hgg�B<̬U(�gܗ^.�do����"��j�1��,�	B�c�5����}$�b:+ž>i;��ߡ��dt�|Φ���P�c1a�����W%�Xu.mG�L"�4��
FܨߏcX�!�`f&H�𿄴_,�}b��5��&�vFl�PY����l�7��Y�����{q��&�����`R�j?���������S4��%!����J�!jMF��`���q�ϯ�Z�-:N��Sth��-Lv�,��j�6w�6�Z��2kF�)�R3�h�"��c���?�C�������9�o6]��Ф��7�Xzr;�aH����!l�+w月�W���]78��q��B�p�=���Bv����
���H�D�6���pS����h`�i��B��T�_�sZC9�s���7�j>�X $���fe/��>U>�����i������3\*�[�MMv8,Oi������t�t7jB�mJ$����ɝ���[Sq=���u�|Ա�oX���)�[	�j��A��P�
Zk����40�:�;��_*�ѽA�<����� &�f�H��(����<U�Y�չ�ޮp�'ƞy�Fd&0l�D��_p�*��`�:z�;�U�^_�`X��s��y��Q�S���R�!.M�R�uLZ3�R�Y|`�;�P�>��`6�V�dx���.�Y#-Sn��j��B�!�Gjf�l��f ��6Y��S�"��2�'u���K����i\�s?^$�sK?��j$�B���(�|[{eS]��"f��aAOyZDٶD!��/Ĺ�Z�r��2�2�7�y��k퓁�3W����B��:bd�٫C�ʠ�0`y�wo@��6q]���5`�u�!-8�:E�U)��3��	�`h�p�G�l � l�[ܒB쪘e����#��ws��fB�����7<�{]^�������W��T�cH�&�����Z�z9�����"K�(�Y�u�;�Ql���
��~�"�m˜f���Uq�_��Wd�`�E���(x*�}�IA�5��]�ev�g-�@�o��x��6��k�
�7�M�+mq����K��ڵo,9�h�?��@���M����#3C�$}��sK�����W�����G˪[ V�.��e��L̓Q���鬃��2�<f�|�i�
���Y�B��qx�y�?aG�'Li��-"��^��'��@ξa������Q��c�tZ���/��Y��I�:w�6ɍ�4�f������՜�� K���c�������z���m���x7�J�G�6�"[�HA�3� 6�F�S �ҩ��=n�V�Nx��o�8 gk�t`�磎�UO��'�I��[c?�T�]��g
�.��v��V�p�|q+���BHj���̙)0˘h}���XRq���Te�[X^�}n4c��[p�Y;ܓ^$����i����D�`*��>�Ѵ�!����X|�^������GLjxa��A(�.ਤ���!�.<��?�U�ܤ�[��c�]9.0����i�Z�������X��`�m`Vސ[Wj&j�����WHvu),�S5��@��N*��>B4�IcY a�m�}X�';'��t!Fs�1�Gb��Ѕ�"g���y��{!E\�:�*�d��S"d�u��5�*<˲�7w��@{�nC�֌����G���z�i�hI*��ا�K��	&�*;�
��`/����M��H�C��xO��ւ����P@��voaL`�����1}:�da5���a:0�kB�����Y<��;(���
A���g���� W�i�r�2��%>EA{=��Z������a�;4��GD�PvHC4��.�&tL糦Nl׉�8�9��K�E��AV��ӵG�,����DW50�t��� ��uې<�Ƈv4_�����,KJ�M��ߒn�y�k7�t#���I�[���R��-/�'$������رE��aly����5P71��4m]��[�D���.k]�a�ߤ|��vB@'a��B���r���]����
�M�ʖi��E=a���?��ܴ���`�L�r9�KE|�.S�MW�p���"t8��c;�ǿRdʅ>u�����.s�:�	ĹA��c����ee���+�#��pxb�@�Lk��tN-:ٯ�e���Xd�e���mD����B<eF�P���`����9E��!L��ֳ�O��j�6�	cY�'�<�*�E&s��xH�d�K��6�In7L�<�X ��ޯSZ������}&bbp� ��~cI�/���/�ek�r%���[v�Ta���H�,~���`R�aW�NU�ֺѝ�ؙt��9�J���c�����v�7��(ER�z2�������Z�9���X/��2����J��g�]�ŧ���hTumɈ��l������+$2�ζ������0�l7s�$1��'��SS�Ŧ��n(�r��T��j&���~�x?�~Z����h@�i��Xc���$��A9t@��@��y$���ϭ������1��=[|p��N�F���'δ�Xq��BG)�N������ю�$��S����A� ����e�K)L}wmX��"@VL���k��5�ݽ�d�F>�兯=X��2kx[x�¥��G�Oz^Zx�r���\f���	Ԛlг�i��7m�����v0&�x	���ny��3<�ՙ��T���6�P<y��n�{t���2��CY<����p�?����jo��by+��7�j�����yĲz4V���`\d��NC���{dL��	��{'4���s�l�v��E,���N�����hJ��?��dڜ��w�-��1������!�F�����# �Γ�N��.�j��,��1�}�?BC�U$u�S�F�\Sň��0~�ؓ\��UK�T_K���?G�$��qiD�"�E��	|�;~��\�ۉ���-�+ć��ڨC���z��W$yƪ�Q`��Ul�"fA�h(���y��Q0gm�ԾҪ|������Bi��!p�n}��p�P]�i|2��-,�/[�	~,�&���D5��Ra��$O@���oJe)�v8��'OV�5μ�z`����k[fGoŊ���J����Ľ���ƪ��SG�����K�rhX�鎟%��=B�_M�H�Jn��.��O;9���T��Y�G$����0)���%������p]�5l	�F|����q�L��82tw��v�:��)��q?�#�WзLʎ�!��4��i�^y?	~���ٮ#)C�v�̌l�o�?��j�
�a3b�m�j$��+��� 6��v��P�c����
7_��M���;�o�
����-��M�x29�B及��S<s���5$ŢA��@�i��@K�>߸C���ؾ�6���_���ܐd�~��:����~����H��U�qAA^�` �ɭ���UfAgE��Ԙ8:5�C;�D�b��3�^aq�(g:�K\�Z\���?��)�~s8�C�Z�5f�d�]8��<���6�ڶ9�`�c���7k��9馰x�Ä�j��}�#u������5��	ym�r�ְ��1����я� �@���LS�x�����`�@�ICk��š���������}�����}B(�N�&Sa�ƏA@���R�	��/������B���[���$*�^ԏZ6�Ȑ�c��f״�':F�c���L)��P-�X�S��N�w�L�B�|�'g,�粑�C��%�E���{r��6y����
-�� ���%�=�����8Η\��^��_��^HFEo+��W��M� ��Įo��Nur@ʠ�ǻWmq��+E�N|�G?�2h��UY�D�L4v@�5�	0���ƎpK�Q�nL,{�ʞʠ'^r,�g*!�~h�3��͖qT�T����Az�`6_��&�@��+,V��6��D_0V¾L�W�ӈ:;o�1�/>tD4�"���>k�#Ȼ�0��T`;�3������ i'��i�m>T濹��r�f�ȑ�b����9?���d�7d�}ǭ^� (�����k���u`[߹�e�E�)�OuW\oC8�;h�Yfk�J�a�Q��4�6&����䡲(�i�Y.�ɒ���֧���p>�8'������x�[^N���~�J�3?���M֯­���^&炠$�ˋl�qk����o�:�%�73F��6�Q~j��b�Q�h��d��z`H�f�G��GB�T�5�<��ZU�g����<fV]{E���7���IM��p�oʂ<�7r�{�*�D�"�ꛁφB��.�Q��rF儳EK˙}�i�j�%��F�UQ�&s�18q��/�2C^�g���з�:�K�OG{J�	e�ƾt���X�m�׌0��\�aV�wУ��n�İ#��f��O�p�50���NgH�l�ۼ��u�s?�zT�!��6�M��l+���&���-LM�I	XWxGtgub���j%�����" �nu�/ՕK.��vPrJ馒�\���VZ� >��
b�6`i�����5������ޥo�f+�薤n'mPqrվ�t�A�΁�~��j�Y�"]|G��ǡ��fkEu����3E٤�F&"]jrX�*�{uk�ˬm��թ��r�2��p *M{3�7?�]2�F뎾c��a���Z��&�
�fJ��l�M��Hi�3aU3��P[���6�9a���q��l#�6�}��)�����x,�!8r�#��������U\�����i���o��l篖}
��Z�_�j姅Q��XݬZW.�22m~RFp���"΄ep7��J%i��޸���=|��ԏ�D�Bds=�� <���ZrMN-�co�+�A���}�
^����$L��gQ�	hO����!�R�j�ڹ���aK�[�h����/�y�Eo۔�lo2�&pWG��Ƹ��v�e��E	��q�[���`>j^�  E�
%J<��oHM@�Z�@��Æ.�"�>���c��%(C��}�B�����K�q����zR��ϫ�J���,x$}ƺ!�Z���y���NR�̚�4��׵$�Q�Ѩ�/>�߸��@�A�c�͵gP+:��D%��3`�	�}*���) g9:�2HS��W�Q��c�SsOz��Ăh�ģ����k�g�$R�lr8�C�7��CZ���rL+��+��:ٿ��t�7�}.���.��~�>�0�	a�����v��9�	�g���T�2�o�U?��q
�G^�l�~mHb���X�oRͅ�rMB/�X9�[z�è�1�9� �s�H^ (2~�+�����������Oxhu�1�g��o��=$:��P�����C�!�E�b�^�񜻟]�����U�@�C#�� gV ��kÄ\t�1�{��~+Bc6�L,��/E�|֘�Z̭-��z:���w�j3f�t�J���*�k$Ι�>"5Vf��h���3o��V3��'���3��F�ݾ�%���7N��2����tVxsهۅ�549�ާ.�D���T�H߶_�r,&4'�lvIBs�D�JI�~��q��f�\�
F��`��lH>} �vaI����[�ℍ�����<
%}9���4(h��&=��=8H*⺾a ��(������;�&A��m��f>6D�NV��pJ��¢��ғ6ٻ�k
@e>������լ�"0�ঔ�����p`�y�ܠ]E�s�04�K���*�g4=���B�ђrt'�fL)֎k��e�kCr[0r�@j��W�`*�vf<��=�t��]7��L� ��t��`ʤ5��"���#���<K�{o,K%��"*Pm3��FCQ�{�Z査x�˯ ����0W�N*�mo��q�H���
��l�w
�;F���#�EG�ć�Ӑ�5Y���!�$�w�$S�S��6D�ܳz�^��D1yŃx7@X{OK�{�H�f���M��GP���]r��I������3A��3�;���G���DN��W����ً�=|x_���z0�s�{>�4끃S<Ύ�Q�3���~(=$N3�8�gH�˙#�f�#D/�.�e�%�d"�1]�������!wp��u6�Qm�o��+���g�#��b���=V��"�����E}K�����X�� ��l:���/�pne+�n�V�d��Vo!w�kS'�9���;��X����@|�{&9�LC�f�RGzΞhbQ/H���eg����Y]Ra�����?���bL5"�Uã[�H��5S�*���sIa�e.o^ڔ��Z�f�ͦ�:�2��m��}v��'w������}�>��%�;NՆ�_���|[/*�dJ\B[	`n)�l��R�{���W_ۉH>�lVC+<��8�?6��AE�d(����+�%.$���1�t瘼E��shejk��T!/:��Qݍ�kۆ]"oq1R���F/K�+�W�Jl���7�A�~ �$	�i��!y���}������כ�c�|x+��+���},M|�wBw�_"bY*c���vb�V�u��uC���nG�u*W��=�7;.+�IvT�1�Ԧ9�T�<��-��!�#L�*��應%7��>B��pu����/5ϱy�������ЦH�_�F�n���\+��<�*��O��Q�����8�^*���e_�ph��-VaI��m�߽Dh�L��`	^S`�������t��-q���^�ſnz��DBFbLb�"\z�;c��Ŝ@E�$�)����l7Q���~�����E 2��t��0�p���;�m�А���e#Kʳ˸��@��Y��/�����<�N�/��}8��C���#obU"{��1'��I_�
#j�xh $�;�d�<-�Ť�ϳ̀��˝�C�Kޜ�����(��kj����\Cz���#-�C�MEk):����K��R�J�:��(nDa��U�B�,�I�x��	�H�66�������(��Hv���Kub5M���9p�8�����%U�YM�MGαe2���B�B���9��Kr�O��I[��l�����=~�mD�d�lZ�\l�,%��4�i���������h�o�E�:,���hZ_
�l��Fӫkx/�����B[�{�x:PAw.��F�	Y&��H���3j+��b�?��13|S�Jt{!�Q��T��6��梙&-����a���gz����!��2�������G8���u�qH+��KM1x��Ե��z��M5��������� 䗒�Î��_�-h��)�������F�QR��;�����e�m�eWY~/��;��@N8��0���#yKC�����D�@"����b�z�I��u\٭=D"x������*/�(��Ҽ=��])	kd����P jQ͚�f�$�g���Q|1MС��%W�c�A���9�J��~�9���b't^4=x��;���G���Þ�ٛRB��#\���y+�K}�7;ZAV# �7C�����F.s��Y�Pғ��#���T(M�&��;:P����qu�a>kHyS�s9lG�i~�C�s��;9�S����4���>g��U�^t��'T�eD4�=��3��=�a >� ��.�_��9��k&�xq,�&W?
�-����ah.ΐ�"�
��lP(�Z��W���d���t�7_����{��U��@�����R]�R�k=���4R��6u�J'z5�M��h
��Og7r��fCރ�!��;Xٖ��M�)|9D����L��m�Jw @�XS6��Q��m�B������]�dbe�p��Ex��<Z��.|f�-��#r����G��2$	!��w^D��X�rVV1��s��u� l����c7�)xN��T�qT)cbMQ��m�>�-����蒻�L��=U��i����6��i%�i�g�f����}.L�J�#��o�kk��Zx����@�+�&�<J���������������'\ͲM�@�E�0��A*�C�}M��Q|��^5������N����*��{;�B'\��A;Y�㰖"�� (	S�?d���]Y�	7���D�ԝ?EM=�UȤ�,��0���p.EE�It�MW�H-_�E�\���p5|CK#�H�Dp��Hg��WC�M/�#Q��wDZa�n�T�󿲫�>�}���/�����>_�
��43;����$�ĿZp�)�I�`���X�� t8N�栻�-�������h����N�����X�TV���f?��|�]��d!4(�6.�p����![�O����2Kډ�WɰA�1�;�w|3�ٞ���Ʋ��sY*��"�B��t�2p 6�Z�,�L#�=�0�ԶL�_:��ÓzNa�) }�0�S�d��m$aG��b�M����8q�z�ߐyf��Y��H	�7d\�����lQ�ȿ�@g��'��ݠ��=�����a���>ō�#ă#r'�=R����1PW���mD�.6r���t:�����G}/o�A?-���g���w��w4{����ƪ�c��\��^o�q�Y����l�o��Ujt;i{u\�a���^�@wA��	�n�sqh(��"M�nM��|�c���;0��k��ZN�O�Z�s��f\'���vĕ��p.|u.�m=`Q��o����L���=OO�c=��k5��re��r5P�N��b�Jr_� k��p&y����[<�u�e(60\@����xFǈ�9ũR��ɋ�~;?��I�f��%���c-^m����6���-1���4K�6΄ɪB�|	iu��%	�47�ʣb���	�	;I�a)�� �����yɨ5��8�DP���Sw���xs�,��)(ihk�iy�,|�$ݧ������}��"��of���ì_��Y����{�_w�#��W��j	�1���Mo�W.%����a/�S��z]���S��։{�|�싁{�D��(,K6A"�^`]p�M��q��z�˦B:�μ�;9A��0j�\8�_s��Ⱦ
>�Y��K2�ւ���^6�$�~0p����~����J�2�P0X���v���b[A,ӟ�?=���#���6y�g�2Rd��S7���(�v}]��:���p$3�
��/P0kOB�C�Y/��vȫ\�yr��<��a��EZ�p5�:�
���,O����l��Z�Im�����L�r���`+�o��-����0��n�}bdM�3��g�@�kH\���pP;�`]�M� ����^�=D��[��x�;ٹ�taɬܔ��y�-'=�N�IK��u��8�L���h3_g�#��u�j��7h�ĝ ����<I{��{;������<]����������f?`,Nl�坲_q���\X�}ԙ�:&�CAX�h���z��!��#�=q3��L�o#�)��� �3>�cX����b��s& ���
� {�x�0�\���R{��$(�����?�, �/o��?RC���I\����#�NY�t��i�}�I�