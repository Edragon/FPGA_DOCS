��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n��<��񩟡@VL�i4}H>��m�/����g.x��/��Ű��	�l*�]��K�Y�D��)��3�]�J�+�a����w�(�� �UD��q��\
�3� ��
�|	I�K���&�Q�Q��8rx��k*��"�X1��|kެ�5��B�,�S!x�����m;L�7J�88˪���)»�vl�hL��6�����,����&���qC|Wd
�!������P�+�<��{2�P�5%i=�[\~�?�N�̂X��k�{����alUK��P��0���DĬ�.t��K;)�E �A�^�y�	�?t�έy��aIc���[=L;�߃��&u�!��~BB#ك��ɔ�*���5g�8��*�C�JXN�@�d~� t�oxg�n�swF���݃��^6!
k��- js3�E�yc�>П�t�n�	~�?��Y���n+����}5�)4p)�QH�	��!���'���͖�~�����]���f�N@�ꂪ��'X)��Mt��z�e�nېe�&Ljꀱ����9@�Y�q��������_9�!5?�x2�J��^�heئ�.�W%W�C1=�C�wd���=���Iq��\�GZ6�sۄk�� �n<�s�_��1��^�!�i���:I9�`��B�ض�x����:��&Wk��1���M�ʌ�-F[W���@n�[WC�FXT�1����ׂ��q��M×;��`%�Ene79����G���O�T<h���a�3�-� 㩆�Fm��YR���:�)d��c^g�d\C9�u��y�\����[�
OS'�:YzŁ�q��v���y �6#iݨ�+p���K[�c���̫���,��Q�� ��#l����,������w�^��:���1��Yk�lAя�rO3��j��4�RR��N��rvZ����m�A=	FMj)e��B��h�k^�4}�.�����"��H�'�T�2�q�1b݂2`n$!
����FhM�m���Y�beM��{	����i�rJX�G{D�O]��c���:nC�;�/���m�3�`g?A�?��B\��vy�7Dpwf`is�Te��V�,b@l��{2�[Q���W����h��'�x���D9�h�Чç���]M~
e3{�F�$����)%y��ܙI̲D�,K��������a��Wy�{�#���8`�Z����T{�$H�F��ʏ�i�?�]��9�z�n	��$��e��hU=i����Jzwy�.�zA�=�����g��9C�%;fh�+��ÿڏ���c�!�,A9^{@U������o��� vΫ�" �k�Dw;)q[�E��WrA9���q���.��("2</��=(��eX���z��,�v;��N5��$���1oAyu����w� ۴j*�p�ȞC�n�#����n�u$��IF4����^e�%�oC�l\��Zۧ�ēx�l���
UWF�f��%<�<���t�+$O��
�2��|F�&���m��u`��J,f�i��D��^��U[�@�����s{�h�a�g�=�2��E���J�'D3�.)�,���1��+�|X�l���M�o� ��鬻�c��d��jz���b~�@�N)3olVm��a'{�)�~ً���@w��Exr+\���#��UgF`7	��7��6R� �q�a: E����2�j��́)Pb��舷�S9����>{���Z�]�
}k��G%�r�y��@Р��%;H�rYP���2�����o�3��6��D4[��@V�"")y�er����Q��AAE�5T!B�~ydb�����'��P����³-�����Ca�B��v�)�2��.]&v�#�"c���)՟/�������Ϧ69_P3�ؔ��5���~̺Ń�hEjB����p���"�A1W��Kt����/v9jN�c���Q7ҋ��
Z���韌�gR�B�X$��U�n�;�gߕ�xv��>�?)����_�3�b\���:�xt Oji� �sɍ�<�mѥ��ȵ�Y�!���2�rn���	�ڋȎ+t���g7׏]�m�kV��-�N�'����F��2<��5����n),f�\8���W}�v�b9�4q޹k�RQ����=�BG���'wc�5��^���g��.vCS��hecǘ�v��,hG~��Ǿ�G��e�rs[���&E��WJ�Tw���|%D��P{a�P1X~��jq]�d�����'�}��ϣ��_mT�LS��5��dw�YRڈ���k��й|㓳	��b��_ YN澳�{�q�����=V�����7ỻ�N��v����ii�]�~��%0T'X�Ϭ7�!E�3�I���Ll'Z,>��r��6�앨�G{��$>��:&}!��<��&���l	E>SZ�qS�gP�&��l �7�T9�w�j�v)	R鍺�G�v����?�e���G'�E���୽��u�gp �f_�������Q|kS��Y�^Bl�/�%�z����^b��p��[�~�W�o�/�ѩ�ɿ�m��(����h�M�M$�@�C<Q�r�Q{����R�@�~����f���r��$��5���s�wLκ�r����H|�t1�U��-�P��9����Ӊ�g�08(�Q��>�"�(�2p%�y�T�������^C��K���,�d�`R`tj���Zoj<���{��{v�b��*���=2��VJ�AB4ʥ����_�.�稴�7ў[�6p��,)���"�ƳB_�+��N�1��c�V��֘�8G�Q�7�$���~�V���?���Ͷ﹬*�������rj���/FD߃�ܥ�2y���wֹbU�����j��z��X��?�K���Gie !�G.�b�];���p�iQh4�r�`�uT�/��R�$��ѓ�Ag��8�蚝~�m�[�V
g����0�u���X� LH_к�1O�a{m9u����Y�b�s&	xC������;gO�N=�θjӮ'G���S0��A}��`�;��u�z�Y�â(�z{H#��x3hP_
�K�X�ڞ�2�ܥy�s�lC��O	x�bt�g��O�a�\S[�9WT��{��^4�:I�X�J.	{�DV:���o��L~p�J���������>W/%�DO���2��u���J���{�����y��> V�fȊ1�I����*��KPV��t(�ům�ͳ�f�]��Ni���Ś	6��~Q���^�8?��:�1��PV�퍲?z��a��Z���[!�3�+��*/{���WZ7�h@eJS3)3�jL���c)�ڠ�cR$o�c�p�]��"�j[N�V��A�MI�\��ޡ�}�ܬ�@ݸU_LC��쁼��~[����ʛf<bd��T���ZAv���o�ߏ%m�Ϯ�I��,�ciu2��["R�A�cؾ8��M%��:c��so_�������7�S��ј�r�e?j�6a[Q�I�,��lw�r|4B =ng��ՙ�3X���K�-F7w��4ؾ�畝�J���_&�����;�U��lu��p��R}i!����JD�-�H��R4�/�.D7`�)4^�5F����1�$XŁȳ��.1d�Fx�I�"�X�6&�D����鿶�F��F��5��O����<�t��Y���4�&hR�+��Aeir���nYm,��`2,f�Q����i�;��N��]�g�_~��R"�I�]�=�ș�����v7���6�ݠ�P�$z����9��&\���	�X�8~|��J����2��#^r'n�4�1�3�<�vSz�?X�T��f`�酞�@��	�^+����k��
6e����f��z�ly�U�w}TbS� ��ζ�yv@W�.�,���dzs���6��$�7(V�~P�ьh��ů�t��|DJ*Q�8��:#�0o؀��ܞ��