��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`nF $ap2JYѤ��6���d`�́ڽ�T��b}
�0?,��n���
�bi���T\+�n������R���� fƽ���J;����H��e�l
��Y��0��"1�L�R��%b���XêD��F�t���,z��{�Dp{C�f��U�}�LX��҅1��I�+�s����$��<f��P��ﬂP�0�I��T ȘA�J������-�&z�q�yX��������7�f[V��}\�u�W���9~�)m蹽V��s���
uG���þ����N8��pd@?����m�<�P�Q���$��2��0	*
t�|o$u����G��S�h�{�ʓ^dԓ�Rus�1�K�/���{V9'����.�2�s�i����A\� k���c��R��Q8�^�=���E
�us�^�G�zNghV�>���hѹ���@����V]��#�n��J�:m�_�2Ћ�P�ŕ���,x�ըWhg�x�'G�/�72�`aj�0������f���b���q��{D��"X�o(��!z50�U�:=�t��.�l���zG��4\spܡ Lq� ��jw���愦��������-V�;�.
�6��w���l�#�DĒA��
w�0�S�>~'�E>hlc�c�pl�N�	���q�1az)�D�乵��aZZV�k
��*$��}���s7�J
�^y�K�������lpP���0�6fo���rh���B�V��m'��;�qVq�9�#�]6?crc����t�,\!��ec{�H�Ÿ�~~���RZ�pj�L�ސ�~t�~�?�_]�t��,\��F�L�viZ�Y2Xe�X��G"�͑��^)�:�Ԁ�Ӵ���^G��!y�[��L���<��]wMkl!�oE����\����"���В�K�c�Yoz�����e�D�!��N������֥!�;(�FN<�����u�t� q �\d�U��q�0V߆�s��E�-��Ms;��w��,P�$��M��!r��#wV��E>ڤ%'��%�N�%%�Q�f���ˍCGE,��T�=��q�6"AXԽbZ!,y>��`�6�z�S��FA��F��$��K+l9<��:�f���j�2]T�\�#���9�6���_%�������a��Kh]S0��i2#���9��C
�*��t݀���ms!��C��ƅ����Z�v��/���,mlצ��{��0�7�}	ݠ�'�(��7�ً��<b���Xl7t�8DI?q�.�ZE�ն��k%������H�	�^!L�8�/�Ff�:�[�z���kMf�m=�Z�/v݌��k}��.�� ��|6p�S+EEe�S��9r���B��o��t��.0+�Y������dJO������.����(�+��K�{=hW�Ëل^�GV�x*7��D����/K���:ikZӔɄ�;��b��1�	�������B�v���� �.�d{�4�u�6��T�Y�G�͛��p�g�2ٜ�8`����ٷQ-�uty��f٭"����,Һ����&a<������N��Un���8,TL��#��������Jl�vGw5�I��m>�I�{��dA9cY����H�pp��3�a���f��',�SQu����M���HZ,�o}��H��d!N!�����������u�Wxm1sɾ��s�:�K�<�CL�Sj��g�Ilvd   �upIP�t/�o�2�3�ř�{w%jJ@��M�mn��q�'ޞA�� p��R����eDV�u��uu��\Xp3+��I�S���8�e`rǆ�X���s��5�%;F��l��������$%A��U61�H4v� A�.�EQ��������
Cv1�n������O��ηq�t��ĪkNy��gc�r-L �pn��A�C�)��t�V�mq'����c���I�:�6�}q�F��jld%���o��-��˵��7�ң(�ޖ�`�ĝ�\���W}�4!b����-d_�a?$+�xͪ�E�ǈ�A��0B��5��f"��x���i��ѩ�������Ters=-�I
7�0K�T�� I�T����=��{��4Ӷ
>$�$�0��x���lL�-"�s�6�w�ò��,Da��W�:i�s��E�
FϨ�����&eJ�-˭SINYW�MK2�>z�
���Nw��Fkc.X���i�5�v�Q����[U�	�2��15(v[D��?�Ѭ�i_����w���a�/�pS%m���z:�I?#����G`}Ŗ/�h.�ˡ���I�H��`�>wa9G�X����q/A/�p+�@A���})M�;|���
�w�n�����]��A�i]qTC>��KUՌ ��A�5�Y�Y�č��Q""r�a�t���rJ��f�N�� db������這k��͠��M/������y��0ԣ��5ƶ��n���s��IDp��nF�ܖx�?���l*�*Nʙ 0���*�ױ2���z��A��ϳ�i�����3���"�i;.��#P+Ѱ�?w��l�����o�ub)Icja�����I5P�lF���T�6J^���_�v7�"ۣ��������$n6�����4Q�����<�b�d��3(mx>h�d�'w��\���9I|r�M1THM�D��H6��o�w�$�_�%�߯P���A͸��h�g�������8<ӕֹ�yV�t(p�}�sK�-\;DV�xɀ!�H���Ļs�w�0�;�D�F�CC�o2@����RPP
�y��}�xiX�ò��5'Ԉ�'I�i�|KB(�&�W��㔕�,�#�KR���J@֖�zrFJ�|�A���<��=_�%�\�&�;��Q�T�=����$���%��
��eL��[�%�M�]TC�%��oz��`(�~���d��f�l���+�q�����8���&�9�d2�(5�-�}�nK��'ߝ��K���d�"��̰�~i
JRJ�f~�U��^k��t��D�<�ס�w\h�~�>0�N�5�ɳ���W�{���m��wٻy���S�׸�G��p�G�1p��M�V?r���2��9zS�ٮJ���x�_<�ƫ�sݶ���c����������e'�I�R�:�+�9-_H�x�]��zc[�HN�'�*���o��k���P�صRX���s��g4�04Չ��H��kC�<����oe(�Y(\W�%��Ac�"���)���M�����'�mFK>�ۛ�Z�D�O���ǉX�Dl����c��v�a�f���I�\8�^E���s9|2��Uo�V3r&u���pg���ԉ,ȣ���je��|s	�bɌÃl�J��-��yB�%=�SB"��&���,�N���+.Ո2^��-J�h�M��Q㲘Nk��s��v�z*�d7��]�1z��=\*�U�f�ws�f��&r���z��s��HxsiS�$��D�x�ZOEKa�����CzȋLLB¶HR+s�H|�3��|E��&Ծ�1�fw�W����	n�L�Y�b��)�ԅ����5\��p�䕇l>(��:��qj�{�z�(�Սg�q-
.|�Ek����X֖���8`=|	�I��o�W�og��X����8�&�%�#�+��]�MW3�[ޠ���#�|�ȧ���{mEN��e����|Fm��&%����N�����*qY9�EE�┮U��VZ�FXF�;���	���zVj4��2�$/�~˺��s�/#A|�N��dO-jʒ�a��X�����J3`�(᭄�n#�2v3ji��?;���δiM罄��0{�V��?}�Du`�O�'V��t��l�I��S��� �� �S %lkX#Cr�ϖ}u��ʈs�WZ󿸝�5�D��ʳ��Ǹ�g-�U�=��`TV�e����a�9?�p��Rx�%c>�h�ۭ:����ސ��	=Ax#�h�3��%کm\�����bY{C
9qCLJ� j�n�WǏR��Q�f����/t����y��A���}8���M��0�5*+TIH�p��I�Ĩ2[�gH
_�B҅06Æ<��B.��Ж�u�Y��}G��'��K��A��9s�rt���K�������Y[����p)���W;�5�_��Jh��"�er��3V,`} qlZ^��}���[u-"w���?��^>& V"_��=�5	�\ �'"�0�K@2���eE�B�3"�[��,x
��}-���t�	�	�w��c����U��glj�8֌�'��� ����M�n���a�v�m�F۟:<�^�A��A�<�T(��цlT)�<X'��[Fc�T�|xL�h�A&e�	�$�dj�0:��PI@(f����V���?CF9v�k��&��00GV�C�h��\[pf�*hoK�������;fx�8&��1��@M`��"x�]0�5qyA�����v��1���me�4�W7��;"�S�6��_x�G<9䉶P짽�#$��)�Y����a����TOob�F9@l͟(��䥥�<�Q��v°{|�f؎�_�7�����~���V��WaW?�>)�ƍZ�C�O��&+���G�K}0�%��H��K�p�%\��]�e��T#xM�s���������_5�e��Oi.��~�X��))!���\�q;ְ������:M0bН�?/2�7#��l6�I��A6�гsň闾�NWW���_Mم#�n�-�'�@C�!�v���HC$��bFP��;�mUg�u��"�r�p5	Ĭ����y*���i��S~H��K�Nn�I6���b<��S �͎�,�Z��%���~$���{��\���۹���U��g���Y�ȫ���`�&,�G����,��� �a$1���l55�{�S���)
�k��� 5���rAy��[_۰���LHb��?�5u?g3M�>+����Ra�����*�����y��G�5�� �`�"�����C�ޮ3Ԃ�j�7/��ڪ]����@~�. yP��h�v��N��f�#l������t�v�&��R��O�=a?=��t�0.S�&��!KF�_I��d���6�@֔ʔ`��-YTۄ�H�S��yr��;��h�+��ȵ,���8��Y��S�(S�9M�i�̚���h��	.����~�"B��x���˧��ԃи�ÿJ���J��5���?��Z8�]v����,������v�4i�˙9��L��������1v�ϸÝ��J��ͫ]�4���;1 ��Ha1|���5���L��#��;�[�j���D�����|d$3O?B�b��$4O���YH��l�dIY
��J�i�y[�i��7+L1�Ƶ���^��8�
{im<Q��#���@雏wZ{���zMo+��	D<��?�zZ2�'�dZ��tz�H��˲��)�n���5(�~?
�t9{���P�GtK�Z-<��FTK�Eqy�ղU|S�ߑu�W͞���`5O m�2�&���1uI���)6Ϩl�߳�`�߄����\i�3P�7��WD+�/����>�Ȍ �:`HC���'��Q�k[-��e�!"jO(���/�y����?��@:�m4.��g6�!���C��x�C����&�����m`{�J<[r ���� ̯kTy�nR_0pn�v�u�����2��7�P�S����+�.l�9 ��t����]�1$����+n���1J9�bh�S6��q�2��lsp�!����p��#O��}��\'z<�Q��jk{H�E2/��_�Yj ���:65���9���RI\��[���]}�m6uY8uY�*�&!t�	�'2-�6����YBxy�31�%r��z8�Ai�.���{�@��K^=���B3����L8�>����ȧ��x���iGW���ea���Hʯm�\��i�� �Z���>�@u.�t���D�O�%��a�בvRzޣ�����c���,���q���iTBH����߭�N�.@�5@�6��y�p+q��6�js�;���K"p詨祔�ţ��������FW�Wb���5Eڞ�P1����u�|��yޞ����#���}.�ֆ^������]���~��H��'�{�YH���J{��}Cu�uçK������^/1�������P�]���	S?��C��� ���E}_0Ϯ2��82�s���JVB	ޟ2�xІ��y��!�B��ȃ!���j��/�a��IP��U�	T����n	��Q�����c�Z���-s0�W���i���0�#>�%q�G�����^5�=mdW${��9ɏ��.��r U*��S��]`�Y�pD��$����(7vv��n1DsE��72����d��_@�Wl��+8*�M^��� KIIE�����xU��{���Z�;FNZ6�X��&�V���gM������J�NPVs ����Տ�/k�֨�G҇����Rp���LOL�򵦙�P�)[�r(� k�u;��1VTFI�������HL��$D1�M��2�0|;;�u�K�$�YQ�<��=�d@�x)��]����Y��+	w:��5t��*K�Ir~��('�s��-��!}���by���̦�
���;(���q�'U.$Ju[��M���n^�y��q3&~��*Vy��%ZP��;<��i�����K��FRC��R�)��^�����J���e�i�ҡ��z�T�;��ܣ�[�tC��7�Q"�__�[���3��n��91�� �禞��GH�bEA��B[��R~g����W�ѯ�/�c��]�@��%I@pk��ʲ+=S|m��1��Ҋ�qe&RiI�(?���q�N}Ft�i^���J����m��)��-�5z�njY��4�h�^�^�Ol%�+��n��jPO�0t����Lr�P�I�^\w���&�qѷ�=���w�M����ڴ�R��]����4e:�OΡXj(�����_��#v��l��'[5t�ג��!�j�8����D�H�H1�,#D��R�����z1/��2�� d�:���M�;W�]��f�q���̖@O��TR��{�
lQQ���z��idkO*ȭb�V�(x�PH��6��C2FU����-,��&ݛwɃ=�c<�w�U�c#���Е�z�>�s���[�1r����`����t$�T�A�?
I���*Q�+���\.��8�S�Q���1�����\�S�&!R6V�/�|�fQ"dxPE�Hz�=��˭��ej�+M�����#�g��[�d�U��1����%�ݙ�҇�"J�vbV
$V��/r�@�w�cn�����ɣ�s3��{R��8�K�ZA �{`��@%��4�-���^6�n�]u�����`	��C1�4�O�ƝV���y�@,PE{�l`c�$T���[��f*/ > �l�a@[P��B{���V�RnQ<|���e=,���/�}
i ����H���mg�I�`���C˷F����������Vm�ý�����gx��/3Q�Úr�丠k�T|ڙ
8����̑�� B��4���=�����<�X��0����z�(�
V8�t���U��T�$8�f"ޟ8{���6�+2I������ozꐆ����_����� y(���T7�֨c�+HFλ�kiu�ġ���cƘ��;���K��0O��=jRȯ�0u�p��
�݊�o|��x�8��v#��2�Z�(��2�k�#
��-����RX��~����~	V
&�Aᛰ�,����9!fB�]��|_�0ƁwE����V�
(��fq!��F¿�N��Z�Z?�N��5h٪<���#zK�t_z�	�7%����2tΧ+�!	ᩱ��J�C	��g�Ax��! %��*�-~�Ĭc��?��H�l�� Co��y��D��'J=C(�>)2TKB�)#��,�jzH(�#��#;�N�x�c9�f?�^�C6f���`q�i��y�`5��D�YIB���>�L8�|�wC�@S5"����@����S-w����#~+��1|�Z�C �����&���PfC�	f<��=�4��E!��rj�%��F(N����uh��C�JāA;�\�B6Q�����t��i-�
PW�K+.���4�.jO�|d���v��xz�
�aa���m<@�L�B��u��@���.Iz��_��I<~F�� U\?�L�����:�gf Ra��)� D8�eB�t��"��[�S��=�Yo�K�K�]�;'�@�^�Ϫ�
5��`�K�uJ8�P�*ʙA�ї�J������HU�*�7؎v�ځ������Qg�Ȱ�/�[0���׾��YK:��6��P���t�W��%~TJ�G�YG�=�Ŕ���C��B]���
.,�����U����L��:���lԂ�8ϗ}a03*kz�14@�u�����շ�M�����<�'���߆��̮�8M��)z�ZL{y�`��p"0��*�a*���l���MQb�WV���օ�*o�r����^@Uc3LB����)$Kx0�&�z�/�,�c*9�C��#����h�d�����zW#���դu���`�f�����S��q��kL�hC��w�Ņ�'(B��9'�V�;��˄��jA9��Yj5�"j0�#xĒs���V�&�|#TD``�F�ް�GsҢ�u;�Ō�����n�?�|[�wքÑ���,�9HX�оX����G��U�P��}����WV�X=e�TF)��@�lp�sϸ��t"� �7#�`��ɖ?.h��N�P�
_���O��\7���I&�f��0�㫘�_�������?�G�TB��!ɲ�tB%.�q^�8U1��4���720 s�|�M�:���)�c�
���o�lh&A9��޶�Nč2u�*��^�HZ�w~C�H��\�����x���/��;�W�B���݈r,�ɕ����-g8�]���W]!Y� h��X�� ��L�u|G���}1����(�F�ڛ|�c>_;���i-�.XD$V�д��f��1W$�%/Qؓ��j����8�����a���M#R�|��Z�4�JV�H�c�ڧdC;o��p	m�)m����ڶE�
o�NM�V�C���7�:g��.�݄+��I�	��=]��!.i������i?-$�*����i@��Y�~��Ʀ+�o ��bF������z�'��62���PK�&w��qH��U��xһ���}��A;�|���F�fXY�����}m�^C�;��Q��=+�	��8������#
,�.OTZ�9Z����DTW�1�z�1�^q�ArL3 ��a�0���z5��p���mk�[6����}�G��B/Ϧ�J�X� n���O�?&��D/g�N���i/RE3\ۍ�i��7��A�&�"W�n-E"ӡ�G�f�Z�8�$�j���S�6Yv���[f$O \�Nu3W����;u�Nx����o�)k-�.���u���E�����;f'O@V��L�T���ވA9l�<e׸A�Ŕ�@�_�Hd�͙pYL��؀�(����{��AzE������;Ӑce�	$��+h�ą������ �v�����h��칬C\5��￭,�-@���lo����[Iˎ��*�Bp���x�j1�g�;��h����w�D&K�!)�!��\.8 7j0�t?�6�C��f�\Y�3�f����U(b��v�=�Vةv(���#���#��Ӯ���a|�O��S&�@�rё������	Fb8�:�+g0��:;��Qָ=7�,�ƌ�@z�VЮ3�_��r}��=-@�h�r$
CQ���k͈d%^�]0���+���l30Ԩ��d���ը��QtO�D�=�@��2����������:E�����4���ș����~�����{�(|z�nQqĉ�����>"�@n2�	d�q˂�q�
���~M�����8�I����.�
K��B�v�,�ߍ�9�=�W �v�T�ԡz��z���j4��_�lN�Q��(N�.*����8u�с6��*~W�W���ݿM'ʾA�j���?���a��w~�G]���~"�O����_=|�J�%çS3*oe	
!�^���{�4nO�K���	 !';HZ�x���������ZwgV����ό��}�Ϯk}�.��V�Pl�-5+ƱB�a[[��P��T�%3O�d	Ԡ�ľ�A�#w0���$�᮹��y��:}�O3�i$��UgއDT��%ec�|�jD����]���$�Tp�m�K�r��uR�Fl�d�������V��5T��q��J[����e&�Ì?�0t�RH +��[���Ï�8Kb`D�E�[:5�TTZ%5Yn��F�M��v�`'�^�w����X6�_I���� ��	̅l������
�,�x̩��	�r��d/q�O���{�������E���cV$��D͉ ����fA鋦���|] nR�;p�qX�Y.vh�e|��輾=�6�GŎ��,�°�PX�^Vۇ��;�������T�k^}�G]�����PV��x��9G�`�Hic+@��<���k�K��L���7��k�%�&.��A��b6V�Q^�~f:��?#|�a��z���I�K-TԳz0i�+�#�)8�˪ZY�س[�v�eh^"E��3�,m���G�h�U��7��l=N�: ��{�5�*~����bY̹{y}q�j���������x���Wv��rq��*��mGK���s;�ff��3q���+�g���7LDk+'	��U�ا3h>(��Yg[x�(��9�l�>H�u�7m>�&\��%�9���OP���7��UZ���q�䈩 -�*d����?I��/��D�)S�J�ԁ��H�S�"	Em5���uS�{��ҩI�1XI�g�V_n�㡦�,N;�Zi�Ԝ ���#��G�ٯɵ:#��m<�mW��������(/�҆4Y��R���>�]F��pbT�O_f
�T3N�`
�=�z�;,�?~+T��k�]/�H�bZ�&���<�
��SÍ��p�&���DB���Wz����ֶ��:㔶ԭ���ӊ���ݓV�	�h\�ˎqq�-!�{R%[h�`�o�>��d$�ۣ"������B�_���
R�� R�!���?7��Wi�6E��VF�;4T�Nwdeuc����
ƍb�I݄��P»C�P�3���z����7V_6Z+�++��Q
�mĒ���D�ɉM�g7�g��`����fP�pNc�&���f�����Vyw;�O����?_{�⩾�n4�ّ�Ex���C�aq� �L}Ƈ ]/Z�k��P�f��/���A��x��o��z���r�f(s0�1꿊��Pu�w���� p-mno\�X���!d�2v��)����D�+�lKz�����鶢�5�tV�.8-~�Q��=�A��uqO�d�9:�v@���}�~��\ZnN�!�q�}È[�M8�0�pj��ї���_V昁�-�Pۭ���=O�u�Y�&b������5��a�_��~ߨ)4�}����g�0Hi�2�+��l33Z��;����B���d�l+g�N�CH}ThTV�G��c�c]1õ n�(��tr�>:%z<�����d(2���O!3PҞ�.7t�������$M�ّЪ��h/�=R���K"��oc����'��l���Pwz�0+�(�?���ɒg���*����X���N a%�,6�d��v表'&��%6���rz��5�»������b`����]��v'@��98�4>��R�yɖ(�SX�f�S����D�d+�py�k�4��gD���I�}Ʊ����5��q�,f j
Jʵu�,V���I�z[v���6��(Ps:����F����}�U	po�59x.�ǁ�ڷ��ƪ#������%���ǟ0��6��L�1 ��>�ӳ���
8�|���+q�-yd�`_�#Vr�O��&jb�|h )C��ڟ��f( ��Ē��ܡ��� ��s+ͳܹ6��'�o������Z
�.����5 ੬�R$d@x3���п���w��J�h��o��X�uЮ�mR1�8s��[G/B�Ԧ��"�o��FXo���|W��4@�=Lt���s�x@�!ʫ"�}���n߲V���	gX[�	�nG����C�򞲿���]�����[+�<�� 
���/�л�Mg��g����k����k��&�h�h�-�*��-Ƚ8��Z�Y5rW~���!&pR[���Qt��1{���75��d�Z�5�U`ڛ��?�_O͐�@�w�dY��,��@O�&i[�	�؉�h%�i�����k��p�~͆::	$:�gO�?��GA��&�~^ �l*Z൦�N~,Ɨ\g>!�-�x��غ��C�� �����J���tGB��,����q���/n��*rD�;VʶXbVb���瞬 ��_.�:�]����6lBnl�P��I�Y�&#M�gm�)2}}͡�|	����%קՐ����Ĵ�.�����!u����Ʋ��b	�ub��.�'ȗ���<���ɻ�?����X�߲�*�U&ex4���;E����[ 2�B�\H����B����O��cP�s�U)���䷣���t�	�ɿ8H8N�3[A�����F	
��{�|�ZoSx�>�����E{$���A��<3#.
��6�����:��~��Dw�����	�4xA��~5�H��U���v\�E�],S<�����C����cP>N��J�-i���\���� U�-V%���q��M��kHS�U��w��5��^��� VH�W=�a�@���bw%	݃Ȼ�����ڥ;7B V��߳B����@�M�0>X�^��D�d� �G�C?�zP�+��	��W��r0�[d��*�lǅ�֌4�μg��$�c����T�׏�E�3s�<�v.=r!E�iXgbb������#�o��?��]�;�(��:(N�X���
5Nڍ�\��o���!�ds��ϘǝM ��;�Yl���+҈�g�z�(U[Y I�J.�ƅ�9�bm���7��]r�(��ur�	�"D��#�� ���e�A����l��X�ㄊS�4%�ھ�:4|u}&��� (k���L>d�� ]ߐ�	��4�$K�Doͨh�!�M��^�'!ϑ�c���/`'t�T 0�'�&x�5��������Cu����Iט��w&A�J.�qJд�\�6.d6b��at�A�ݝp�H�FqMYq���KLZD7%N댓� ��&T.r�2Xj�Z�3o�T�%�5CQ���x�Y�&[4�w��������8���(�]�]���
R��b��Nn���ue���󹲡�+*���*�/Q:v�M�N�lA�;�[�Rhj�kA\�2��d	���u�0߁�ý��5�q�\�G�4�>�� �:-��!�bn;�÷A�gR&���\R�'V�Q�ixj��2:�?�~
(�^�܀�A�eʥJr��7Q��XH�Vh�fLG~ɻ��F�T��R���h :Wm��'��14$�Cs�S/�hW,�.��KB���'�+�Pa�I�OE��2��$�1�+�>�&/��S�zN��1���������9Pe�aë�~o�0Y F��'�gH����SEߗ3>�V��*	aJ��� ���.ӝN�G��	��CL�*c�<��H"S�u�\^|X�4�����0BwU�{��z��X��I���Be}l��~$�ù1vpts���h���j��{���q�9I�Q���;�j�F��0��Q�l�=��tl%[�_6������B�]|��)���y�:�q�f�L��F��:�}T]߂fB��ɠ̧aG
�I2 Rt�{����/B�J�y&���v��{f5��"���wT�d
F��l�<�`��X�a����沒Ď���]��d�!��>��|)SS����Y���d��	C�}� ��={׹3��4¡���dZ�ڄ���t��h
dbg:�Rh���CÐ�'���Y�W^g�h��6�=�E�@D�/�
f\��2���U�5�����/}�v�q�D��RK�n�>�����:n���"\ �
���3�7(�𳱫�:��LfrJʡ7qx_�V��9�o��W^hx�r3՝�%�tlQi]��Do������A�u���c��Ν���e !R�p �����C꙱������6����҇��]ш(/�s�g�B��T[_���-�[r	"z|�w�đϊ���I���:}������ �]�B�	�Q���];/;��a!D0��w<(����m������U�#y�p�'I��y��8}����m�K�-�3��. ��1�.�lL�_T��}�28;t���e�a����Z�_���a�w��H����a�|j��ƵWJ4�,kא��D�fz!�͂�-_����X/���\";V��*��֜!�A(����:H�����	�����N�R�mf�t_��\M~����p*v��q�(@-��ː��p� �\����bk7�U)��%$�p�[�����M5��vE��vU�GѦ����T���V�Ms��4�6�����ZOx~��2��q¿�6XV����DFK0������g�/ԍ�+�8$��4ra��M%H�ُ߆i`��n����5��[�ȡ��We�Q�1� � ��BJNP�{Wq��G�;X&Ɯ��r|N0��W��?F�O�N�ۺ�bos�~��6D)���	�,���M��xrK��	a�Q����BL��ڒ!67���9A�:m�b}<�ʃ#�dݒ����|[ ����ҍ��,`����^aj
��qǄe��`߁�.> ����1�gВ4���j�1���l8�w���������v>�m�70��$|�:(~\��]�e�q�M,&�2���R?�S�"x�q^�ED`�����\�!ɶ��?�
��my(Pl߀�e���3��$,�^7p@�4h��ۃ��+��e�)���p�F�#KU�S��)���U������C����l�,��~��Z�z��Z#MB��ԫyy���f۸}�ǟQh�{�Iv d��-��pR����/��� <)�����Q��:/U��w$=�k�ub	���K�<Foݶ �^�q2G�^�����(u0�I�D����7R#9n�[A:O�t���,��P�Q��'�;ӿB�%e���[�'��zֽ�E'FPH�l�DpK��9z�
��&�X=�-�L1u߉�y�%.���?�F/�.�$�tޣ�}�]��?�G�/��h�-�յ�#�
G�$n��6�1�K�0Q������}�aUH��{_�4���l ��J��z�8��y���{�&�r������}�����2hCR��1���w~�M)�)���_%�(��䚞Q�k"����ٽ	a9/����j�e{S� A%��w#����x�͢��"�	W��vQ��R�������"�����ޜ����b�֥�QS�a�_�ɯ�U�^F�9�h�I�Ov���꼋B:�o��Yn����o���P��0��CM=�Y�����_q��N5���_���4V��=���sd�P�&������AM��@H=d��]���Ц�;�F΁U�<�&�6�y�.�7������ғŀߊ�Ka��[�8�\���i����|���P���5�*:�@�`��3�ꔄ���Z���Ah�v�
Jn�c���:��WT�/��ap�_��+�=�$��k�ʕ��.�ԣ х!��F|��gޣ�^lL�b���v��YK�o4�����&�_Y�"w�,��:o���Kw�a ��bb�[�|K���o��a �جu�����h��h1�W�A�u��P�����@%T��<�u#��N8C�ZL�k�C�"�n�/��(�uO��3Oס/��JeJÜ�I_�H�{c�M=	[ �5Ls0�|xNs2?�^-��ƏP=9�^3���r���"��Aw�3"bI�LQ�TC�Fȅ�ܨ�l�P�dr��`cm���s�����;:x��Db��v�h�΅~������qF����+�T�m��e+*5S&uϜ��[�­ˢ5�/�|�,�v�`7&�~pzZL���7}O��5qM�q��!ꘈ�n�8�yee���R��&6р7�G�|�׀*���"�b��{7�F.SSux�������7K�@�(��Y�zNgW����9,�9��"a�mX�TjIa�Y�4���po��=o1���L,����p7��*{d������j�:�s���9�V��Qj6����H-=�TM�vRj2	OR�U�ަ��i�ݪ�
Q�<s�J��ʂ��C[p�o-�oQ+Y�nS���܃��Qmn��<s�a��bW������Ջ��;��h��7w�*<h�_��H�q�Jrj�0c�s�i����j�&�;}I��ߎ߭��	:I��OR�#@Kl���z��1a%|&��V~rή:�� $z̒`��t�x*�Vg��p�t���[�ܢ��2�+&f�Q�G�qy=~_D�� ��^�]��K�epS���?c�Gͱ�BNf�Pi��6B��Uc�����$��ʳ�lx;�v'	]���̀᣾�b�rg� �uU�:
l��1��*M���� �d��:X�E�CCdA��.��!���rFJ�¦�Y��i�x���-{�窧w� �=��C�$X��=܁���E< ��c�|ǖ�DFWc����4I?����eJk���$��7�+�)�e!�ݡ��I�%I�2�6
0"���Ag�A�C��j�;���E|�u���츱	�J�tq�cH���]6�V@F���� ��ɼ:����<�ߝW'��>B��}PM�LҴI�6�n���m1Ɂ����Wֳf�s`��o��sD��O��ͼ�OrVAb�g�ת�p��@FYK+@�f^�G/�C���r{-ӫ����;c�yqA}��ԥ�ܥ�-��Y��L�5kg#
�f
��+=��љp� ����լ���Ay�ׯ4X/��tYMy	4i4J#b(g�7��`�qY3�͆� �*ca�R�/��VW�,a�m9���H�5�ȸB,���i[�󪞀���̌��l���r�I��8VR|d�A�WG2%y���2�b���vvu��p�4$�)iH���$I�>�;�頮*ݗw��4�W�*h,�$��s����r�<�p�������G-�O�}�L"��0D�D��ᜉX�G�%�Q�=�K�����%���'I�~~?���
�j�7�d��y��*wd�m�&����:U����R���s@P��y��"<�z�z�Y/D�ar�M���'��v�'�S��{z{(^zҧ5 β�Ǹ�8��49L*�([�Ȫ�y�:��aN���s��9��D8�kpT�4����ޗ�ў�m;�G%Ӱp�1 S1�R.Y���˚L�I�3��@֯c�yJOw)��8x#�Ց��3?� ��/%k���u��b�`�MT�d2��v;�bk˪x�Ve \'Q��56�qyU������6繥���U�R������qb2UK�
����3VI�� �뗒���պa2O�7l�+���\t�y���-����(���TJe��egJ�NJ��R	])�'$j��epl�\b�*`z�#u��W�/�z�z&��Cl�Ү��)�cЅ�K�M^��YS�Lhg:�%Vtm��g���� I�^u豬�ҖF�`�������pR�0��i�OV��#��y��dI�/�R���ڌ�",El_W_HQ�ORѧq�ϻ�"X��Ё9X�;$.$D��x�����V��۪2p
�ỹ�e ��O��I�6kܘA�f��"q��є�	@�ht=��=v�4�OR>�R���R�]eP_�F; �2;t\�rQ�*i28��p�1���z/t;HWC�1ptv�=�Ι�a��FzE���T�߼�8���E��J��|?e�CR���.~���r|����4Ԥ|��X�*X-�Lo6>?����� ��t�/�}�
�w!
����'#��K�'���1���
��k�a���x���o����vH0z V��߂> ��z�8�j��i���'Y�&���>�y!]WU�
��@F�}n���R�|Y]z�a��4����^\C[��TH?��6�m ��ο�G�X��:�X�Mh:D7|'��q���C=�Z��9�@I���v�
ߌ��6����4 ̱�E��X�<�>�}��� ��7���4��*�A�NM@Zhu��l�KE}<�l�
դ�	�������w�(���p2���D�r7&�~�}�=®��q���+�&��[���`���I��ESU��yS!qÄ<��U����?�x�$M�Q�%C��l�E|�3[� �ĊT��͜T���8��i[zS�Ȩ�Nԓ����{�wD���g�w�d�2 ��ٹ�ۓ��꺍���߽�$.)�X|����Z`�����"�@VPY����T}w��k��n�Y�|�Bg59+vI�恇:�ڳ�i�e�X�t�pL	���!��O��A���Ex�ّ�<b~��=ۥ����-�n�fĆ�P��m8�&:eͅ�����8�	����S+;�� �9��i������?�噼�c-96����	٬�mb�x�K���KVeWi���+Ԗ��-7Uo�$16���i�zJ���U<���F�E�?-vc8�5����X�=Rm��Ybh���[ȫw�U^�j�uZ�M�ܾ����떛J��At�~�&�v��24yw���à���<���A������fn�`�rR�x���s����d��><�sj'�@h�-Y�'�υX�o����$���C��¤�h���*E��[}���	N@�< �ڦ�e�>`��
�?�hjh��eĄ���qz��_r;�)�Eol#i�S�Oyxڗ�6�3���33��b��W����A	T�h@��G���+��t43�Uͺ�$ӫ�3CSEq�RKg�e���8�ҩ�!�=%Xr쮥�Ŝ�{�N��O���'`4r]�*���T)ҽ�?����d0��l��Nu�Bf�� �1��!�I����.�m��Y"���A�t��P+���� y���N���ߏux=O� �nX��j��"?�l�I�ֵ5N�����zuՍHҩ�(R�I���I�pA�䅋��Y+4�b�L���>76�🄽u����Yٮt�D֥��"���\Gdt�������o�b���{ؐNU��	��0+�_�L�o�!B;�H�F���B��Рw�rVg����F��ڵ>�&+�F�	���������, ��A]}�Xf��T;
�@+���ߴ
�~�m"�>�� �)�����[�\��z(��I�ޅ�� �"�LW��q�𿾄�7ٰh�a��-`������ގutح��͢Zj���l_����#�u��Z�O�R:D��M9j}4y�h��)���������"�u�@\� ��'��-�J��is�V��@�l���p$#��C�J�W����������#�$Q��e�?l�s*8�Z�I�<����2������D���C��(Ȅ=@�3}�̈�,ܽ+�btuҿ��v�F��h>�7�4uh�Q|`!��P�Az�^��;�k�L���~B E�xy9�����	g�<�xÉ0�|���קSi�'m3���_�PG�4)&�cX�L�?YS�hQ|��D������Uq���;H��=�dI,��]�{�{uM6l�u�Z=l�C�a�@�9{4�ε`/�<r�5�;�T��GVs/�R���������m+�[9�ȓo^y��=���M5JA
��7z��8�e��A�N6N�b�h\��]Y6n�B*��	�fӻk���I���x_��+��TC���?�_��:v9�
��%���2��.�&����_��u��o��H,���5�\YXh4r�(-s,ʠ�8Yc?dMp��C��[��ҿ�U�} c��x���z�Y=U��ҟ�6�D�	��i���3���$|+���dO��/��9�\C�ՠ���o�5���c�u`"4E"k��C��|[�V|=�����O�$K)̈D����!6;��_~��$=�TG�
�L�e�b��lLwU��,k�6��}�E+�0��8�V|�hor3�]�������|�YlT���*���ߛS�>!;��b?㟉�k��ݦ��K��1$2���&� WJY���F���E�,�@%�{�h���䂞�&�&Μu�p]M�!��E5�����k���JV"Z�h^o���
����}���Β;]�&@�Q�Q$,/'���+�h�੩�:����(��ӱ�`D9���Glv�g��UR��a0I")LY��z̍�2�d؍B��q�A�NRw���E�7gW���Ӥ��-�ֹ����A+a�Œ���Ύ��-@1zKU���8�B,\���/�{4����!\���H�^|�*sU�s����Y�R����Mk�\�����yZ	��O��Ҭ�(�s�r�����61�I�86�Ыmu�K.�ޣ������3j�'ۗ0��ZcR+�]4��*���Ȩ�_�2h���1b���n��8;�3Q�Bѵ�/x˷ɭ,������kn8p����pv
u
m��쇣-K��������"N7,�wGť`r<�MM@a���Fa_��������r��2�,��>@��k���i���^�H]R�e����+���'���4B�ۡ*�NKys�<��K<��XC�@�O7ƙm��_��8�0�G ���d���~����G�N�*<���q+xP��>�[��7���y�?�hi��B��~!d5[3���5x߱-J1�tp谯iEY�������o� ��A�JC�|�`fa�*}	���Y69���9N�y�����w��?6����i��9ڥ3��d8jk9Ԥ�e��
X�#��A�^%�q< $��:5�׆&���a宨&:~XD¿�3����7��Ԫb �^����d".�-b�P��z��*��lY+�*]S6/��O���:��t!f�F�Od�q#1'��=�*Cx��U@08���|T������`����8[ȗ�z�k���N>���ώ�ـ|v�+�/�4D���]dJ�q$ [=9���Q�*"����@���/�	��;�I��QZ�2j�t-i�d����%I��l���ESA����tߏ�#]�oy�(Zざ�ن�IfD�ԊÄ�:���ԟD�%*�+BJ7��i�d�����h��zX����^WD/�M,��.�Gq0��?UR�@O��A%�Ȑ��7I��X��������v�b}���-���Ny�@98H�3�Yw��8A�mioJ�O�~.�xf�E_�9�Ja��1�u��������b��@ic�v��:S��[΢;��V���(ѐ�Y+0s-�C;�%�]97���s���\*G1_���1(c�?��[�M�E%��Wr�Ea��؂����pU{�L.����rv+`O$��d���h�]qE�t����R(!���"}��EAzCD�xtם�;�d�(*;�G�=�ش)��� �B���Ǎ�-瓥N� `m����D�%���Z�;�ZTB�(����;�_[�����d!&�9Nsb� �����t�Q��(���<�pi�ni� 9[H��M�l���h�ޓI��pR�F�."#��>X$�o�)���p���s$e�/�>�Y#�AuyA��Xsٰ�������Hyة�"�=&�;��e� 0��ʺ�YX��{W.zu]V*��7��ׁ/�����o���)�/K|��šH&HI��d�Zp")@j�h������{>����X���0^X���&��������g^��<�-!�)t��T�.\���8��M�'��R��Q��j�	nl��s�rp�.�~"y�1�+��#��J>-��	�b��vW:)�?�l{s���;a��9	����5�5�o���d���5V��Ya��S��f���6��}�DX��cc��G�Vk���XԸ-���͋V� F̵�?��r�v���E7���䟠r����$j�^֫w���2�W�?e�~��V[��+9��ԥS��>] �� (BC�����dw���	�\^��ǽ�^]�nG�h�U�Id*�j7ʖJ�x���JE/4BAKkMh	����f�d��tiי�}5��Yoo�F�5+�:z�[��ZM�X���8!I����QX0>��/T�>�� �O���)I��i�9o90Q��ձ��m�&D� g������<����Ւu]r:��n@�黮R�B\�N9��	���e��q�IM�-(h�B�l��l	�Ot���a�?��'���8��+���UB���*>��k�Ñ`/����R����މ�{�[s�Ѩ-T%LҶ�9�
� �n@R�X�5�(>z�ֻ(dw������v�9jw���Y��*g�/$�wI塔犸��ڗ�1G!vb����+�U댰@��K��o.�q�ȺĈ�A~�ӛ��律��Bk"�}�oU9d����q��p����#�������q<ǒ�]91��(�Ii��j8�I�Sp&m��Ԍl۠z�\�ʜ� )�����+����g	������72���W>v��)/�+��)�eK����c��S���l����h��슇 !ddIOo�Y�5|CN/)��V�_\o�e	�0?���c}c���_�qD��.~	�v��Y�o^b{cW������\��]@���0������ӈH�du����~�����[�ԐR���=�̒1Z��B0�;v�-ۧ�y�,;���v����m��ނ�(��m��t����Wmi�ZbU(y��Z��+�x�k5�$�*z�۩X���G�+zïL��U��'`qR@�I�'�v�p;!�!F����D��s���F�D�����d1�~�X���f�!�� (1Bf��|gj��y�
���^X���
�.��$8�z)�1$J�0���g��)�07�}K�o���)��?$�^�'��!t$����7?�wu�������v�ޜ�(�;�%Ec[CŮ���X��K���\у*�Xf����D<�N�ۚ��[*M�>�'�y2��7��r8��2�����B.!�g#"��#�}@ӷ�8N�A���ȃ�	����=F{��T��jg�̓�Q��;r����\�_�rLQ,� t�Ed�w�3��| z������g�O�$�;Ζ����\3���������x5�}X����Y�(t�!C����F]�C��
䩧�f��v�~j,�=�gid��J᭺���fI��s�w��Nq�D��/n�q�n>����	�ab����`��B���5�i�Ș�E�t��39����\��U�$�I�J<��tf�ӈ��c�v����q�H�K��B���w)��{�'֣Iu�&ܰ�ם��zbQ�V%$W̦��4�ۤ��w�ңç�NQ�R"Ĵș�����h��܉�l��<��t���h�@����5��Q��� q�УYeS����92�6I6*���Z��y֎z�'-/a�X��X��	�-�!Z����}$b`���;Nە��ntJ��6̏������%�v�Tҗ�m����/gZ7��]=.$�ur :����mj�U��-���_���+ұ�
�����X�l��ʈ�!q#�*Iq��f7z�W��:gNl/��O˷��$[��/�à��|�c(t��F%~�]Rxc����6/�˫}l>ԧ�3�����$��@<��
���:�z�\����}=��B����I2�f�I@��D`�����48�nk�ڋ覲˱l�4j��S��k��˻�J�hi��h���R���ps�)���xoM��'��F�6B��x��TV��NJ���P9ܠU�z��k訁I�(Ch�#K�#J��+r�b�0�M`�����9mT%�;��M�d�H_���k5鴁sZ�����1���G�L�ra��e���p�J�f����r���\.\~!"u����F�N�9r<�S.`����*+��%�@�����Ύ�}�Э����y�5����m�����F�y�d���#��
}�D� �"'�K&� 0a���f׀�<��m[7�$h+)ȫ��4���$M�M��{���@�y)-�n��m[�)�SS�X�Y�G�p��Ǆʹ����h�.g�R��d���N�C��>;��4�T�~8Xe�ՙ���}�;�+�3����	�\�Jݕ�������o���얪:wjǙ��l����[؉VPk�x
��l��?� ��+�ٚ�����uo�֢%?l丸D�I�6k��#��{�����7�Rm�	���h��P粝��d�uƏ�F�d,�t���̶�C��M��|G���68�z�.��F�S����.<�����>P�2U���1ߧi�9��_�|w��h����J�W�0_/�'--VS�][�y�X��I"ӄ��&�+������d�B�d-j�z�U͢��33���c5��~v3�SX���vM$j�z�����C�;r��06�ZP��Ns�ɵ�l2�o��0�����K�LZk�����cF�뛝�`���c�{"4��kde�K���n����_B�'�2F�5��������[����e����o�w��u1��~��G"6�$k�0>��4��kt�6�����g�H�K]�$晶K�Й��}`)�S��s�O#/E�Ýs���<��=]<�&�D'o�