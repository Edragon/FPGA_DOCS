library verilog;
use verilog.vl_types.all;
entity pll_ram_tb is
end pll_ram_tb;
