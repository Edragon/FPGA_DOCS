library verilog;
use verilog.vl_types.all;
entity altera_device_families is
end altera_device_families;
