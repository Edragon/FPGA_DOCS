��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`nR�D�&�|����ꏮ�f���oX��A�b��(>��ށꄱ�>_
_��Z&��r���8�'@h�T�=���6��K�`I#��Ǹb8��b���.C�ȼ��tl��X~sƪ��0�Ԏ1&n���׈�&�{��m���Kj.3ғĚ\�{�STK�C��?�H�W=�t��im1�r,;�P������ҋ�G�tc}�:�b����HK&��4���/}"1s�Ѡ	4�NV�&J�	�Ƥ�yg���n&�D4���lf��N�V�k��7�0/�M�_L����9S���h�9�;���l0}$���<��_�4����(/;"����B��0C�E��bY��;�����h!����btp�%:� �n܋���8�ˉ�O�֓��B�6�Wȟ`��p��� ԓ�FM�@���T
M�X�b�>��g��X��]k�c,���T8V��Up9�������f�qh���i�c�^��醋�����C���o>���x-��A/�����uJA�c֝!)���k��˴�z�*�:�79y(�M>���+�vD��	O0��ҿݺ�w{�G���sI�:�.G��W>�!W���	��3/ ���TRr���~��
v�++B���G��
��t�6�ĳ��V~ tN?c��[ʵU}*0?s�-\N�ª�?��,@\q��,]j}?�+S�v8/$ˋr�f��I>�t��M��+�m�"'�k�!c����N3�`�u{Ί�q�t����2t?N��{?@��`����.������wB���"� 洲�`��v�F�K��z�3��l�\�<C<�UZ�O��C�.���T�Moj�0��R8�$�KA�n�8��Xh�:|n�V�@{=/�4���_Tr�)��(+�B�<�O�dL3t>ۆ\|�U���I�B;ؐ��Q��$�7ΥʳR+"p��wD�=�����P"%�@s]�R�]U�%��u3Ƨ�����x0@+�~[��L���t�.�H��/jL��B�*댩Lv�vO=~8���6d���o���-Ԣ& ��q`#;r�OO��;Ś�!�,o:i�hT�ZL�*#������ȶ�l:/$��:v6U�^|�@^is�#�-�'�5�$[dN_��U ���è6Ce�S�"|�	z�P6A�z�b����8/a:G9ZD�sF6i6���������y��pWJ�wч(���������Q�ROL�<��(��~A?;��׿�A�ta��4A��b��JH�X�b�Sm٬8�\�A]�7;�N��R�E�Q5��1bN1�H�"�Lp�����^��rj拑��z3��=�)�N^�/�����_J\�������6�l�G�Y��#��A��'��Np����o�#����#��4���l{�1��0������h.������J�c�/�|-�<G</��q��#�yD���H��W���K_�F�B	���.B�1�ǆs�O��Q��scf__�"PǄ�AF�4{~�w�?s	����-�n�RZ��H ������ee�fB���*��Z���\ ��xė'}��__����=��{��ӚD���~`�NY��BJU�^��P���������a���Q7ɹ`�f`�T׾��2�]�N�`G�!�>���3%b5�/��>gUM���2\mť�j��9{ar��z*�'M˩�o���잷���ԏ��^*��C�Kꓔ�"���||_��V�ͬ��vn�S��T��`��F�� ���ko��7�S%�x��!%S��9�e�����y.�31��#�3)�%
��0t>/�ͮ��)m�U��mWs���_O�J�����䐂L��O�S Q��uW�2�)V��J�i%�� ��{�ƌ5th��ę� �?����������D"˿����A;:maXʐ��c���&�m;�BV@�LH����Ο	|��1f����F�,	��5P`sh�Q��l5�O�wr��F%�
��Y�ѻHg��l��a�� �k��*�}I�&�z��`����8u�z��r��`����(�5(�r����
���t�r��Yۗf6�d�B䑏��ۨ�5�1���4ob���I��]�F'�����/#8�Ǝ8�@�akW� �|���~�QWQ(�Ra�۽�>U|�\�@؟��º�)NfS���)��@���:>Y���Ǣ2���=��Y&�%O��a��#��襵�s;�����vO��X�NVp�E2d`mg~�*�K=��֐.ͲOۊ��ؚ�lrE����\����5�z~��� e�+�x���5�g��C��L*�H	tWgp�b䅭cEE$�;�g9���y��ܭ�.eb?���dW�����CS�]*�y�h��_�&�1�}0���uD%_B��h)�~=ȯP6ƹ�mD��8q�:�(��^aD(�q�U�3�7^r܀%"����/�#Llp^��~{�}eJQfS�j��'�Y?MѬΌ�|2��CY� ��t5��=�����~[ӱP����5d;��L-=;�i4��e���s3�����[� KfYM�B'�#�r�]����|���j7�*Ⱦ�<��T�"�->������4Q��v�'�{<��$��Qw���=�t��b����b��'s���cœ�X��H'�@Q*��/� 9�����b��;;����n+\{�߄�>\�9fWW	����.�ڮ���`��[�X&��N�Г�������UMi� �w��?&Z���j��Q���{�u7>z
��S����k�R2�����;Mf��,T�_�Ѵmy)�BqI�xnGL���	4 ���Q�SY# �����'UvkcY=�w�����O�B�.�=ޑ6c�}��Bg�1n$�?��4(�P�$��D"���4�֢��u<
Q')vԫ[�Zx�t0�.�,I����"���:`>َ1���&��W��:���7tAPBM�������Ή��S�K,�/.���-c��I�X%ѐ�����1�M�����l���1�&�V���}q�)6�(�r@�ofVT��Z�U��K��L��QFƇ����SEv<���1����Ŕ�q��D�M�1$CH���5���v,0З�a�n�(�#+x����w��Cpe����*�m�X���]N�B�r��I�\�++���e��x�@�����%�K��_�)(�/8�M�euҽ8[�Հ8+��	�m�y�,'l�q��%���۞�����_J��yY���m/<b�rz���|ӣ<XWH^h��!(����u윿Z�E�n�:N�3�]4�@=�Y��E<����,#��qŋ�g���ז�h+0X�������^b��l�7��"�R��;����X��43YiB8[r��	�G!��~��x�o�ʛ�M&&Wl�+��%Y�-���QK2�ʮ�������B����]��Z�tʰO.�v��*@�X`�W�_�J�s�'x�&�+BA��ݯ��,3]��S(y�U�O�t���q�����314R`��YC~�?�޿e��2�:O��p�ڄ��'��|����wNsǥjm��6撓r�o�!��5�Ho��tDpdͫ��<��Xۿ���9�\���@|K���X������h4������<x�.Kx[�T�=
�4]��Y]oD	����\�7Y0���f�4�nq<�X�4p��.�C����&�22Ώ�,�؜�b��8t�Ǖ'�`�a~ �K(�2�{񠢉t�]ىΞ,��o�Qa�7ǲ.��C%���$��{>��C�O�V�'�?@ܓ��G���Ƈ��K�Bd�WW+h�NZ9�����'��5z;<a�S���X�����|@%���&~V3av��49���~��:[)U�x�~�0i4�&~��
�O�$����moS#i�f!�`�ٯHpX|��/:d�.� �����1�R�]W�In��G��1'��\Y�xRX�i~�!�Q�u�7*'�F���Y�a��M��Z�;}`���X^]Q�	g���%��ݽ�-��g���;�bAq�{����-��𥻗�|�8��SF�lf
��V8R�G G�+��p����;�L���Bj��b����ʟnJr����Z����rj@��JX6%�\S<��F���Q�n�@f-R*�R����=�p�p�/���}k ���&�k������m�YJ�[�6�(�Ll�zn��t������X��^YAX.=,��S�"-���2p�N��<�9*�V��L����f����*�� �H�l�1���O
�_`S�4[4=��F�"j���`��4�/��	wÆ�*�r�B�����ΏW����Ĩ�(|><s��b�|$���d�ۺ^|p2fO�M���:y/Ƨr+�!�yn�r�Z]�N���u
��?�L�0d1��4.���ӫ������>�t���F�=��l.P��6wp���j���/[a���um^A�c3��W�O?���yd�����	K�!k�Y	��s|l�T�J��9|��
�`ί5�� �i��o�|�'Q�uH�8������nkw`��&iGPS,�\,%�l��Զ��:YmŒ�T������Mp^?P��v�>��H0,oْP\�J�У�E_F�	u��gEW�6kK�L94�K�����������:��l>�Xc-u�ĐK3@��Ŧ������,5��I�P2��l��wb���߹���j����wKA��X�cr�5��d�����j�?�	~E^y����yC���V�o�Ђ���4��6���d�|�nt&���˫-���d��{`���!�\��Ջ� ��3M�B�����E���~�ذ�8,�WV�JM�e���3���:w������ R���vd�Ym��M�Cy��oR�_
Q���9�T�mck���c�b/��,
1#���#C�ab��
j@��3.ǟ?�!Ǧ�s��B�	�E��ֻ�p�?�����)W��1�2û��qs����ϣϩt��-y��c��+�n�|�S�{�pI�ww� ENؙP�>e��3�U��7�����̩��8�ww}�:�#701k�h/�5a��p�۰d�n��rߢ�o$�v��+��������>�*A������`B&���eB�
dvV��e�ăZ��_�Dl6GyEd��۟!vzwt�[	Վ�K��"�bs�k�F즚14�Q;d�d9��W�j���#!X�v�Bs�,E~k3ە;ujU�vPeɌa2P��Յ'�L�N���0�w��H�W0Ո�I� ���O�{w���=�DxW�����U��0�K�0,X.���w�U��|&��}.B��H ֟��*�����:��h������{sVeN���'n�V��y��+�o7�:������}S�D����X�9��R�;]�G��*���P�B�#��ߛ��u���a��T�xno>������s}��
�<nl��b�J.�T����<�3�$�j���K��O�
���T�h\�|�-(��y�,4�6%c��2� ���Ss�yd̑�9��M6�J��̙���x��=HV����Ľ݋hE�� �,!-4�zb�L��c�WB�0^�^2$���/d��V��(e�G��'�M7ڣ�t&�Ә�`��h}�č#�	sE;t�a�މqb�$�L:�7+���Wߝ�?�$%�`H��[�j���o�g�1�\,ȇ`�݅��[�rvA�yx�7:��a9@���EI���m+
+��Wq���`�x�S^��C�v�۴��Ԟg����ʫ��wBd��}dU�7�H�ml��r��W�v�h�y^�޳��}D-Ge�S�V�􉁍�m@n���;nD\��f>���XlU� ��Գ ����8�O����u�9Mb,����вi%�k�ُ;'��eǴyh� ��r���튇�h��,^��a�=R>mfcLSz:	��A�8ǆ�I�8�	��֏~`�iA5yښu]ѭ(�
����z�]�eۮK���*��h3�� }������}R�g5�����x�<�:��|ƀq�ڗ��y+�AH��|s9 8cm�7��c�)�0�\q ��a�c%PR�K[�=�mTH�g٘���<�e���W�Ef��	K:�u�^��	xnt�wթo"��1��陼�&l�a����m:M�{ ����9���C8��������Z�2�Y~�+�08�[��F��,�QP�0h���t��ǔ�f����K����^���}3�+*�kO4�g�op]y��s�o&�`��&^�t�e��H%FXA�k�@��:�I!�)�ܩ]~��D,�ك�#q���@�ϫ�kt\{�IF�<��"=�f.����}�C��P��m�q�
cŌ���5֍0�)��oΈIn�FJ���5��[���D��t����8P{ �&»�A{;���z����5g>��ݕ��s'vB��q���j5��|c�Ɍ�M`�A|6Bc�5�`T�X�Ҍ�KҘ��2�O���l�bw-�WG��ɜ�ޅ�ۑ�
��a��{�`Έs�^G���y�Nj:�����yX��}j���q��l���YR�E���>3O�����!�p�E��ke�#l���5(��y�︾��9mzu�����kئ�
��`3<wG�s���O8�&�`�'=�z��X;MҴ.w�q�$�}g$����HM��5E�X��)}"-���a�TlHj�R�2ϋ�z&t[�C�;��e�J,�L#�v�Z�F�׳aZ�c��1u�yO��R�c��ÔBf�`�3���zX��M��a�ߑ{���Zj�nC)�'L9I��@_J�B@�xc`'���LK��%7�	�b4%��{d�l�S�h�T"��|X��O�"���KR��6Et�<n ��%�#����<K�AS�Ep"��L{����U>�����a�T~a9m�?�`�����<,<ܻ�ݜ�j��8��Χ)m�;�<u�m�r��7j)�vIy��}6Y����| 2��NE��9�zY	9��
_��q8Y�O��ÕNO�!Q-�4���� �u�=�H�.:=R�/h$��.|4 x�Hj�$��hC�l~�O�� �e�^.h��)��:d�p�����}6no�n|˭UH�KZq4Q��)�B!K�`+�j��q
G ����]`#���S���Dj����[���O�/Ga�o�ҹ��n���=�?�J�Z%ћ�+�����3��J��	򂢹�Aн�����7�A�`.�����)ԯv��	ׄ������)��a��H���`#с�Y�l�?��$�!��
U�,�� ��a����?���4t��݋l���,�Z�ۑ1BH;��N��.�SQl8e L~Qjs�L�h�*g�|���V�� �b7�W0��`_���7��ڷ�dl����:��	A/�?�-g*E�'��Vz��)y.�Wt%�c��ﻪ^�T?p�O��~�ƫ���WZ��3���]v����\_�3��Ȕ��.N�81W�m]��v
  314�цV)QAꐰ�S�cH���w�.�A��0��6��A��񏅭��T���/0�Cg#�����Ύ�?;�WG8OG���-������-' �\ƪ��Y��]|:�+K�)#���5G�y-�F
_���<>ʼ��rQ��vF�4p�RM�U8�sq9��f��_���/1e�O��Yh����6���V�4՟jL���7}�+q�,�O�D<����%�x ���U?�
ܿ���;0������HЛ��H����Y:p�p&�g_g!Ŧ������@~��v�澱@13��	6���'��9}�1i���^7��#��k���h����v��t���
�T�{Xܹ�~�=���M���Wk�<��9h��wB/ 8m�3;]�e��{�^�و���#"k_�����rȩ�Hs��� �x "?tg(�04�Dz��"mϗ���~ʂ��j���Po:�"�'. s	��}]u��#Z�r�@��`��2�����P�'�Pc��! �t���a��?@��N��r�vg�`R�ϥyqƚyG3�NA�ߴ�g�������<�<�3��z� &ǯ�M5J��,�!���"&S�;�R�4��5C��$`Ug&�WiZ��G��O|R�/���:n�-��
oN`
Y�I��0ڠ��ƈ�9�����`MO�(���sf��)k�l��,��~�Ć����3g�Gm���A��ėAP}96\�~���s�A���d ip�a��ЋRy�J�$U�5�MY����/xB��t����JŪ�]�6o�H>_��]'(�N	5����ŷr=���_�ǁ:�t`Jj����J��xP�D�.ͭ�5��C#ԍ1N|�L&d�'$Z�8
�B�#ȉ5Jn��2��&4��}��}��|���YzR2���$���a���Hʔ�	�:��a��H�Ez����Bi�~��:d���a�h�@���m����-<�왩���\�A�'�r�gk`9
Yjo��,wf��U�aɡ7�Z��=>��qOm�7 ����b���r:��[��5�n%/�ʅ�e-b��ݣU��vZt�����C�p����`a���{�n��L�^֒�����������=	�v�q��0)M�YC��=�(����~ƽ��
Ռ�]��������!�;d��7~|��D���q*�x�6�n�=�	����;ϒmt�X�JԤ���}���c�f�}A�]��Bp+C�	�2p��]�"�u��^�{.��!�yEo����kH������9w;K{P�A�J�#�*{+z�l�������<xuW�����K�jO�����˦W�y؊��gy0�S���~�����	"�벾��k����"���~Cg����D�54�����pF�z��J]�LƾDׇ�A��p������S�ֲ���N�N*���5="<��E���''A�	~l��.�Hz�b1�4y����W7��kQ((I�<��3���">��y�B�;:p�ӆ�T|R�o�wCU]�T�ZI��ƺE�ޙr֒���g�)0H�S�h�s����z>w�,
3�2A��JA�äY�$S������(�E�Av�n�TC��~�k�b���o�T�=�p���](3�k�*��d*%�8�xdm���%C��b�~�ur>=6���pc�欜y�^훫���a��1,&��.ݲ�C��U��^&��6�T�C{`�'X�W�p��~U#e�X�4���$#���/�-�k�f���A9�I��շ��_�:�Ԩ�a}���4)`8�Z�����uF���gF=�����pa!?�ꀛ��6����S�]�>�=IE�Bn�5��	s'(�i�%t
��RA5�qpU=�/�iL��p���:CD]����Ds��#�Dx:J;]�a��S@�}d���\5no��i
�'qbw�����o�1��rQ�}��Gx�Ķ���T�@�Ӹ��;���@~�W�z�OV ����73M��W�j�p
���bT:�Ji��<lG�h@vbS����c�XP��,�����_���=�Q���S�6
�X�bg����D3�X>�K9q n��j@��rj�5�*�ȼ�ܒM���Ey��U��}�j�Ix�����M�� �JJŲGm��g���>�vٽ|�*g�5���Q�K���oF����H�8�Ov�}؁^3��K��_���G���<����.@�x����Tw���<H��R�A>J��RqTG��׬��� -�NT�(��0�_��0V�?��� ��
w?����ޢ�����wB�O��h^asypg������K�v�z��Z�O���1�R ������=����2�Sg���r��R���쮋�����'tP�˨A�#9W�F��"��gŔJ�q�"��q�7�>�އrFbܲh��wq��x��ס�F�+�V()J����6WH�ÅU�0�*nA��/<-�*�l�Ie�Թ<m��xy��N�.�ߊu(�\��-K�i@O��b�c��v89n<b�i�@`��X��lpݭ�%�m����J[���ՀQ�����
��|�b�\�0he�ֱ�,�'�%���:UWEY��>�v��^/�����u��b:h踜���;�ȿeeI7�`�q��s�mL�yY+�豈��P]_HN.]yfJ�� 02�<	J8GB��;j�&�P^%E�^�Bn�JB�×�t�&@�QUk㱬�ȏ��f��c�B>���li�i�-�T������g�a���d�ͺ���8�ku����`j�7i�ʒL�����n�>V#ID���E���E�K�'���`9;�JB��E�J6�R�Ϣ����+�у���[����<W��XH��Jݠ���j٫�����`Q��zԺ���=�O�J��^�߅����^#���壎�����V&�B��꜈BY[){߂dCZ�~�,�U=R,ޜ/ �%�R�ȶ�_�5��`%}��8Y��b�.������A��G���*�@�2���!�����yQ_��^e�_n�q?^��7Z��+�����|g��%랸G~,ղ�i���V�B�^���6�t
gk�]������nl��6F-zz�d�De�D�e����i�3�Q=�
����|J򿅆1x5p�:�\ᚶ�����D���]�=X���9��f�-�A���Z�6ac� ���]H*4��%GP��ۃ5.�0���3C{s�پ�yg,{&�h/��E��e���I���Xp��O><P�׈���Lj֭���n��76��� �ۣ�@lu�s�I�����?H����_Ғy��c�<k�R֋�w�o���ϡ��u��魧m�h�0:�2�C�4P6�y�#�X=�`��8����u����.U������Ko)[��Q0�k�pkz�FdY�'?p�߇���e�o���H<�vW(�i�Қ&G"^+��(��gh1�)I!�yӑPTM�^A��K	�'.ݠ@a��L놚j|�0?�zY%'��O5B���F�Lw�;�.杹xea\M��g�G��O�ɓX����#tﻼ
Y�Z���gT�.��ʴld�l�OD�T�����6DZ"���.;�VB�`o3��ڞB��u�̭����E8�9;9c��za�5�(eD�$�,)j~+7�"Bl��l��O���;|	WƱ�K�ǁ�JSK���9��.����D��@O�^�ZP)\��^�6��쵹ל��y��wۀ���,�pCcY�Q�/jSv����%�l�@nǞO7���0���?�N�H#������*�HV�)4�	�Ӥ??ݘ���ќ��W����B���c�~����K����z%uw|= ��+T()-��#��|���c����(ȡ܊w��8���.0�8p�UP���6��D��Uh�穾 ��d�KM�y+�19����%�P~��
��E��o����1�>�p�4+�cPŜ����Kr*;֬xjX��Q���S�оQ�J}E��{�q�c1(e�参kl-�8OJ�Z�H�c	�Z�F���E�wso!h�DZ7CaO�C����o+�S�j��eϥ�Ph�OL�V쀴^�Ս��!2M�[�(܎�#_t��i-[�h�M���&O0���U�$w�T-˿(r쒘�X���)3��+��u,d��~����8}�4�躘~Ӂ�w�⺑:S21��NƠ4!i�&4�vC�_7��u�!S�H��a��JeJ�����208C�&Tҧ��9羺3�0��?a�iܨ�M��� ܏��Gw �m�������E�oR���h9�WfOMExh�\W�TK���)�>C�=�+r㢪g�d,"D�ћ��a��BRu�JC�X
M�P��9L���ݝ3{.�,���Ϲy"`	D�*@5C{�N11�f�}�*F���
���߬��n-�gC��xV�v�]�?���;b���<�n�E���B��/侧�2��Ӟ«B�'���������Y��6WpTj��uO�s�U"��$U:;O"�A��S@�XH?��Ɣ���c���|7/#u�����JU9A0\"�6�T�[dI|� 7�������L�id_'�īSרQ��@�+ч>�}Ъ��$b|���{k%�{�6�n���ka�� 3�Gz�O��W����}͋BD�t�����t~����w��O�4^����Wl3!N�n�Ժ�0�۱�Y�c4�M$A�w��lm|�$3�d^�;��� pl9]����GQ25�Mu[d)�\�#�Y��V�F?3�(w>$����R��]��S�e�έןV��m֎|&��(�I��)��� �H$�?�[���$Ng<*'u��2��z�}Q"����_����ҙ4�tx�%G���:h�Up�CلRHy���2��#O�%x���!u�ٱ�*ab��9�E�8�9O'6�}�"�������nZF���m�����-�2#�B��l$��% � �3�{1R~!��XLz+��
qeM-�"�rM?�~��M>*hq��,¿#SM]*���{�܀4~djR1VȈ������G۰��!�!����!{ZE*7�*?�B�w����--������I�GZ��g����X]o��r���Nu(�&��|�F�Ax�I��/���|N�R�GuN����Gm7oa&�UmY���t�.ƖC[�����zJ)r�c��p�]܈�kR[��c�>�}�^2�)��9����n����7Τ��|C�L�L�t�d��>�*��0oKR�8ę6�WXw�FM�V�rd������&R}�-`Fˆ�M��l*ڋ�d�Zls�G$��mS�(�y����Bz2k.q���`3t����.�sUa/��^�_�YA�ܛK��r$<zd�] ϛ�/�������RxD��n�5Es�� �,X��jQQ6��H�7�����Ӧ�eR�vB�<�t�>���n&;�#h���u��l;q%?W�|�o��=O���.��,��j9x��������fO�M41O��L{��ʸ&ol�� ��%�p��X���ˋ��+�$�$pv���.�5�jj�E�a�=��զ���r|$ ��� ��g��S���F�=�`sI���-�[R��H�߳�ãIq�|���� �e�~� �~��XkFኋ���%������|�!�'�HOH���7�� �ѫ�7xo�������CՐ�)c��Ի���dQ[���KL�0��G�>~~�J��H7�~���4KzG�N��;��wD�wx�P�ط1YS��t�3̌����<a$e �fSzd��r����%J�8Jt�!�ʐ�_���s�ў��vS]H�w�g�rNY#B�Z3�O�L�~��LL.>d1�k��;{�+����/=��.(U�#��oA��F/5��6#����c-/�O���~(x���2(��}��e�t�&�Ke��/��`Tp�A�ɢ3����1�8�O�D�:Ns�l�?�~$����b�lo� T���g��N(�w�J�������tJ⽣f�3���!5���9A�}��w��l���]�	�E�ٺ�ņ$@���t�Lx�Ґ͵�e���]S_[MQN��h��Aѭ!G����YO���j��bh\���~�TK�2}��'��Ҙs�T;�G=ح�够Qx��.�WaQ�!:��J�e���}����a�8F���f
锁<�Y��N��p��l�$T�K�?r���2��;ڟK�	\j`~]7i��8�A�	b����?�H)N3%n|���涺���t]� `��%��eTDH���m���Y[\�as�͒���K�1�Rr7��_�F�lW�v���*��2�r��+��\86��1���"ު�����A�\�OorzE*V�4KU��@bb0I�X{E��ߚ	�dk�(���%HM��@w9g`�I�b
���0γ���� @��p�S^�97��Ǧ�������_=�=���#KٴɅ"���
H@�8;Zɯ��gF5	���A����zB�9�-G��wl�s�S]��U���gk�_n���$��<�G^�>��Q?�HE�Fi�3w<e(�7��p�u�������d�\"��\��Y��M�~�]\�iItH���F�"��E����]_�P�ޯ�bQ�S�h|�R��������W�r&�Փ%�\�9h�
�,��0ZV�G ���;��;m*���Fp��c�.f5n��������y�CL�fcYT s[��Z��V�u����Y0m�Z�j�	t��t�����ʌ���V�g�cQ��,8b�U���DT��9/�h�B����,Ln4�}d����٠�
�ۆg6"5�k�|����yi 2l�>`��L�b����O'�^�|��XNƚL��ռ_Zy>۲:yQ�L[�R���I��Z�D8^�ҩ{NKwl�OLK����)��>}�k/Z?���gs��s� �s�ǂ@a>%z�:�tg`�|����v$��3���$�C`�ڴT�@��\F6PۏG��gOT�i���3E����2j��CV.�$����XS�PH?�2�7�ߊ�|-��=��_�6h��'2;�����
���PZewM����}.W������Έ��zF��z8'V���g� I���"h'^`��ZC�E�	#-twᐔ2X�d�5H21�/��̫ �;��g�1��41 ��2C���aBi6�5�CּP�C����)�2N�+�p��:���X�ژƾ#lzuٲf�Pƙ5ewA		`5�s���E*\��V���˳��V��L����"&W��������X��f�������}���ƨo3ñ��|�/Z�_q��ֽe�;�1�؆��(w,tS�vS�³2Ll���^R���#&l�l�%����'��ei��[-OG���*�øR�˔J����f�Mz�h�X0�"��:�ŜE)ۙW�z��� �v�;v8$Đ��گ��W*u�,���l})��,C����g$F��vR�b�*Jw�|�� L"���Y�Hz��.K�p�0N��}��)KdK�bx@_Y�7p��]��!�c�Y}l�\
f���>�~�˕��f��V٨H8l�V1�2�X¢��#�	�]�N]�-�Ga4�t���`
6a=������1�U\���Y3��:��0���h#�����V�p����N�c�.ɵé%��@��� �P��j����?D�Y� ����6@�D��Q���Ct�6���{u(q��mU�����g���zއM6�+���<$В�w�3\�*Wa@�хpßl�1����&��L�{���4�D�%6������A��ӭ*-팮��~jܓ"7{Q�,sK�e�΍������(:?d��ɒ_�>��T����h~&�^m�ZŞ��o�f5��O�� TѤ�[�;CbR4Xp]ePv' ��z�ƂVƌ�k�2��8�1;���DwO(-e ���ڙ�w�]��y����9�ה������R{�﫭V����&��=�P�Gz�8٤�޶��s�*b���[K��\����o[Χ
�g#�	�Dq
F���ߖ!I���8�1�3��;p���fF���W�\%*�$�2�� ���@M�̃�0R$�>��/�f'N.!#��Œ���f�n��PB[2)
e=�p�5�0��Dzb`�ĥ��*۶�:�y�w���%Ĥk�)�$SŶ�V��CWzf[S��Js�;�e_]P��9���{��]t��!^:I����,
��
u}ҟت?4l�Θ�R��-@|���H�u֚���r�2��G���=!W�`jӓU��K������|�N,;�I�,)��Y�ܢ.�#Q�E�*�7N%W+�����֢טo�dRu��&��v���u���������Me��۴XJ�w�|؂�[�P�Mi�?��`	�.�0Cs�p5=@ c��r�{��|-K� �s�� A9S���Çt���Wd�v��p�)5��E�ϐƯԞ'*8c-C�;�f+xQ�"�l޶"���5��U�N���b�+'"o 	ԒT�?Lb�	�	��c��uiv�ui��U�.(C|)s�E���E�?Hn9C�T�.��1�ͫ��ۮ��r��2��j`MPj]����α^����MZ&(䪧.��:I�rz��C�������ٹ�r��02z6KS���!hL�O�uF��B0���v$�!�-��{JW#�H*�=��oq�K��9����e�������,X?+
�~PN1��{�a����� �@7��G�qz�{\������n��Dy��g�`CO]����ޭ���P�X�
�~��rd'�]Z{G��2>�f埳��� �S	���_�1PG�R�7Z�*�>��Zi�!<L-)/S����I2 ��Sm� p�0���EHj�!{�a�z�A��J/��,�&1�8�No��Q$�q�����ԃ�j�'�$�	dM�Ww3,��;:#?��X��e�p��0/�&��Т�W{�j���/�r�b2	[2CU�8�@4*�m#9ק�8��Դ���-��k̴q>pa_��	�k���#�t:=R���k�ot��GR�d�)	��z�&��˾v��x4J[l���I�l]��u�@1�&��
��t��v��$��+	+����5x�!`t����۫<1��s`. ��5�ȻCn;��
~�IPB,F�1q|���N���C[Q�T����:���Д�0q_�����Nѽ��tc֐F���K����! ���`��vӷ����˅J����]EW�j%�
#���UKS>�����s$�����®+7�  ��6 ���P����.-����D/cМ�g샃���1��%��W�d����;� ޥ�����h:N��{~۝�T&W:�J�����XX[�~d��|U[b��	JB�~25q�Z��j�V�dNY�Ӯ��X��3BE��o7Wq�n��<�Z�b�X��4U�T�_�k(8������Y0
�]�����-+�m.��:bhVy�Ɩn�}$~\��!��3�DWl��� �P�y���;*س<�L"h�1/}7�C�T�Q�O1�/��x��^��pZIW���h�D����@��M�x�E�3
�0ɑi{�ɑ�rD��� ����K.�\�)���P�p��Ip�S+s�]w]R�_�pt§��`�����8|��x*Y��3:I����=��$1R�z
5
=�|x��ܴ�U˴0��"̡`���,=�2+#.F[T,���}�4�P��3�7���� P�E������h ����
�B^JB��K*24�
[�m�zW�[rctK�e!�/.q� ��?V�pF��L��\�e�����з� *ns��\Ft��d���Q�5@ �_��s6��{�Cڢ���pZLӒ@�^�f ����O�;[:p(�|�XS6���*�jEʠ���D�VDk�A8f��T�P��ex����"Lk�A��Ú�=[ɢ��%��@`+�����0\��Spf|Cj�2�v�W��R87<¨��%.��麭�7*����P�DQ��}>����=�Oju�]�	F�~i�ty~i��GJ�[h5�3p4� �o�,T�'J���t<�|�P��u����,E�t�P���#U��jU�j����:�O��#8r��G�l�9B�W������,�����	A��-vz>l��������>]HG�\F6623��^��/��\j��b�����ݪN1�޹�a;�XV��4�6�j��i��~���G�����bjA$�A�R�x��;�ͦ�XT���@h��lA�?D�?u*,%�ߍT���MI=D �/!40��V�`2�����&�]
�aty��"!�:W���o��į���8�wM�;�>V��cvN ~��Ymiff7;
�˕���U�����0�M6���_�%&�k�6� *���$��*`���沜��
)�øx)_�u��i��<��K�*�]�\�S�-~dP֥`4�w�(+
�x��Ti/��`o/�����c+ۿ��R'���+�b-�D�3�>���,;��l�u�pԡ�����0g�c>xoI˾���c�؁�ӗf�WUPSw�Q<c~���z�rk���+8�y��N/M�J.��&�Ax(A1�2���+J>Q��/�?�PGJ�D��|1i�_4I����S��Vܝ�a��K��1��W��!r;A�MW��N�	2ُ;B��,+�6���3���XR�k�K�(㼮D1���?��)��C?Z�砘���~r )'���?Wpl��G�w����, &i��i&��W����:�}@ �L_"�"TX��d��MK����l4F�$Z���wD�����%r���B@./�l����'[l��"���z���=倱hlJ.��7T/�{�����EZ�Y�w��h��9�����K������/���1¬=gB_~�:�S�\��R���W�/L�J�O��m�hh�"�`6�$2���_l��^|J��\&�zMJ�d�]�Y��R`CA�����{gX	�A?�t�B�V{=\@�;O%��E�	�YXwi��T�E�7�bp���}#���k[�cH;���#�PպԿ�D�����G���3�u�c����üq�ߑÿ߄x���r��~�X;��Z9��Bǔ�N� b+�H��R$���?3���L@�e�>b�>p��ж8��'�>�#=�g�i�n	Q�� K3�d�X���m��T�[}>#�"�)��L�={�q����Q����%�=7�<҂:�f=zV�<8Ъ5D��_7R�h)mk����Y�� O�B��.�.����u0R�Ei,�X���7,��ok#
����Z��m�ܝ��q���H؀�"2H0��ȊB�~��3����O����kZ%�Ύ���>W�N(�x\�;~-p��d#�u���j��7��&���=�}X��SoU��i��P9oˆ�.��[mZ��-��(�ve��6�����_���M���^͡�AI�9S.|�N�k '�\;!�4�̽��P�4R)-*Xs( �+p������y��Q���t,�����m��BcH�ky��ld3@0��=����4��~����YM����o7K
�{�s]���L�
�B��KRZh7hKL#r����6G��¢��x��*D�i����W?z��'�?��ؔl��Gx���!ͥDg:g�*�Sb4��]�EdD1Awv�>��ڢQ(OD'F����T7 �E!�u����{�}줰5U��[���G�,�c�P�Yl�������m-����g>M�LJ�� r�J��׊��d�.b����	�����D�!)�8�����\�`��Q�%5�V�.�����9����j��R�����H���/�/Eū�`זl���0�t�`��Mϴ/d�;!"X�.	xy��:uL(�'�y���Z�r~�v������LU�N�}��ř�v{��^��Z���˯����T3����!��]#w�fM���0�#�́������5�@�:���%�p��1=�Cѿ�O�H�4��ݞ|U<�N�7n8��3_�p2[��L��W�hd���K�	�� ��X����3����v�p��㻼��ѡU�&� �B��V��`����4s@��3rN���+�|*��O�ʱ��v�u�ŒD/�5��ѽP跇A�of�kӀ�X �	�f8+`��:G���~+��!zmB�����6yñe��᝽6�p#��P�7��`}��3��f�,3 a�#�� y}Sa�_Áx`_���.���s��KZ뻳6����jtyZ ��_P���/\p�*��m�aHV��#��DQ6Su��M���Wzō_$�|Lb�S0�3��Q�d�[~c<$�зDB��L_�f�?曻oGb������* _8� M��e���+�#���Ȕ�n4`�hnJ�� �,��͞и�|�qG9����6��#�	!��{2��u��8GQ���(�� �!�ՋrO>��V1�oY�$��Zc%���h�K��5�U���� ��H��`�*��θ1��)o���`C��rB���B�0QP+�8���e�C2H�j�k��k:���{f��Δ�����۲�N�d�F���;<���81�_f�Sjd��]� �ֲO�پ���n�b�����g�ƅ1�n)R+۠��ZK��N�� {h�T�a����X����+G-�<9�d��[���o���
Ɂ��+kP�g]��EM(�KK(�s�'��=ĹԴ��w
��py	A��{�G���\-��{���6��*����i�Q\��΀J<Pu=�LP�`��rp{.$(�tܶ�������٠k��{�:t��V	Xm������gC;Uo�H�u;�� �XW|{���ATS��bi��ꮀ�Λ]�7�X䰹�B��� �޲ZR�z�;�������'�O�1����Ǹ^��{v�..��]u;���Nn��ʣ�1���g$�bz��o.ڡ`�0>�����%D�qXA��$g�yD]���In��2j�W�e��G�X��)�A "v��_�{n[2.+Y�b� O*�5��j�S�Z�""t&H��#����-�;j��*f����#SN5��� ��Lls����**��W�F�22��Y;�FN(k��ļ�3���D�
zssM^���7���+E��U��?��o$[��;���K
[J�g�*K���܊��� #Dp��/�H�̢cʎt�!�7ۣ�g�BH��5�P6�w�߭���D~GO	�"�)�����PS��Do��4g���촷����β���
��J�3�=�;���!*������I��nk�����S�O~={��.��W�)-/X�	2�|�fP���}FN{�I�$R�a?`-�"_/�T�����G� ��BC�u&si	%R��OK� ����s��g͖c��ji�6-:@~��gC�ؕ�`6˂G�r��/W�V�����EюX)Ca�m��5Se���B'Sҧ��.H�0�y����G�V6�:��
�������mI�Q��Q�6M�06���K�]�� 3��2M.�E�\�l�%�CC����1� �K�P�B���Q6���.�,�_�}�G)x���]UГx'Hk0��o8�x�(�\%O;��db���Q��#Z��kD).�"\���uI���M�RA�%S��®rd���3z����^�V�i��9�xX�[��HC�?���|tRt���O�F������!И+�͛Pz}h�W���'Pl=���oB�#�������M�ޕB�{��PU0�,aQ2*�]�J��� 	G����q�Nϕ�a�����	�k��i/��l��&^��&�p�ݬ��ȩ���ei,�C�ӧlpV�x��v#e'^4-���֐�|�:U�0���I��B�Q�SȠf-k߷�Mߐ���L���	�RYDUp*0�Y�����r%~\?�QLZ��IF�����Y�x���"�=�z��w���7=~� �
��x��]b�/)л^$���%�U4'Td�F%�c�9����h-�M�_�T,Cpʓ���x��ty3����6-�!=M~��'��f��r	d�Ɯ�:�*�,36�µ ��m?@ڒ�|3a���v�{F��X��}UË~o3<bO`���*2M����ˆ<�[��H��N[�!ʣ��IN�9OK�[�/Y~%�L�G,Q����L��=B�F��d��m�b�!d+�8��0)���Z$u\�����]�7�P�g�M�*��,���{h�>;��g?"��N%R������N´�x2A뚸A��C��D�4��|~�w�	�I�t)�T��#똩�\��iQb�sn�q� %V
�+]B��s~�h|�~oU�2�Ü�rƗ�������w����}��,Kv�H;������C>�
�q������6�N�h�;��.��}%?��Jc������B*|��
z�����jj�c�R��һ.�Ew��"��h$�&�(���Q|��e�S���#pxy�Mc�ԩWds�sv�弾�x�+��f���zPmb�H�?������4x���JJ��*��I�yP"%��1�t�h�7����mc��
]�er���I����ՐW�	����h������M�@C�z���@)1)�?�L��z����s�XE�Wgt������_n��������G�mq�4��e&��A��R)�Ugd:���m<��[:�<؜�΢b��l$�[}����Å�@�Z��T� ���vh�)�֝����{����i���\�T,��1�ˏ��=hljC�2h,�(�3F�� ��!�\�^�$�u��Wꢾ�986��mDd7�张P�tUh(�"a%Q���C>����)$�Ϭk���]�\,�c�c��|G�2P�иfM���Y�`����f��1,[H~�<�o���~��ߒmY���8�T�]�
�3j�ӵ*b7P�ÖT������9n�Ȧ���"z̆��� M'ª{?�E��]2Ro�iW��]0£�<\�h��耸�����W������Ϩ��oU�5�x�dɢ�_�I{�L�D�oi�ǽ�Pn���}i�#w����y$��P:���w~�5%4nt�� hGn1�m_��><��zY*�0/I�L�TVΔ�~k=��q�*/˥~Gϖu ]T^��7��_YƸz���3�{rR��"(���I�9qP��ĨǠ�ʕ
�ݹ�8�yX+�����kS�%ey]�\�{��_��?�H_z���Bjp�H<#�9a�܈!���T!5@3��,�����4�P�'�����}�w�(ǽM�5h���a ��+�J�ƃ��
Y�W������l�'�Y2oؑ�o(%��>JvϾz�hH(s�i|$��Ԣ��O\�7ee�M��Xm��F� r���̔����H*���ߤ�ElP�s�-A�h��V4��]?
���ӖD�@�,�^b��'�E2=�k˙� �����_�IE>7��9š�zX.Cp��]�-���Y�AS��E�+��.c�4
��rg���HX/&��)��h��� [վ7Ԁ�z�|��ƍ�dȊ��lټ̈́�>,�m�M�5��}-.�9:Q;0Z������G�s"�;�~i,�"?m�����Y�#��+�jb�e16z�(%6���>�[iL߽���b���X;Tã0�'�s����,�~&y�|�Q�?@/S���ݜYֽ�� A˛��7y�㥩Bwf`�Djx��R�35�o� ����h�C�%yN2ՠ��]�.�Z
�����#�4�*S�YaK��^�*�Z� #��`|5r~(�L$gUc�����+ ��e߸ ag�p;T�rd��i�c��Gq�c4a��:�O�G9�Y]��R�5���>�E�*�2\��fy���f�n��ծ1�v��>ۛ��z��J�l�@G}+�]��v�]m�� ����U�8�E����$��/�5?-jBs2���+s觤!i�F�҃����V�%��${�z�,m�Kcj�D0�����qŚn��[�]�G��^�C�߲�^-�\+;��@�T��TJ����[��<g��B(��5��:��#^��is�K�aK�Я��4��Ӓ�䓘@=��,r	]��I0���5- Z���=�����7<6��p��[��1
��36ݶp�j�q�k,T��3�e��>N �t2s.�K�ߗC�N,\\�Vqx�-��OxFʉc̦��a�H�����fJEc�R]��Y�Y��B
5��	�y���'Zv;�SI3ؐQ���X둸��(Q�
��Xa�K����L��H��p��Zf)��e@5&���"�Jf4�����a}#aBSL�k#+���w�d��O�4������������޿KG���[�r�G�cv[R�4�4ƿr*~5	)�'�4�s�rP�Tv�e��\�p��h�N�g�m��J�a4�3�:�4�~��H�a�P�˹�;w��y���.��$㻬�S��	�^�,\���|�0��UH�����o�L�,L©j2lY[�q�C���cO��a��]"�п�t�G�w���+�c� ���j�ڃ�K���E����6�!�@��|�����#ǫ�;��D�}��n�Iݻ��X��_�P�V��5�\�_$�A��=�%lcɝ�ÞG�.�j��A���xa�yݺ���)�ӹ��U��z���s��}��kѨ8�wT�ߢ�@��t޶R�V��^
6�[ۨȇ���y�h¼��@�N)��B��U+�Ia���,����.Қ���7�ر����\ZW�������릔�U�D@����E�@�,��¤K�.��e�[�8����@H�����C5s�<�X���%n���vd`�c�����Ru�V�=��(�C��3��`�2��|�����B�UE�m��*k���W~?���k�Z�M7csK�]$���V��F�"ݧ�n�Ni��j�6�eiñ�)�9�[,��<��a�X����u���I�i������4(cշ��&o%��N_Y<{ 3r3�����1�O�*�j�q�6ʒQ�L� �lh��/�-{U,%�s�!�5��čC��#���\b�02��߄p��7�ɪl>Dh0{��" �c4du���F���̂iH����Y+z��as32�������ݾN�ϼ�S��^6����W�1E�6��my��ڷ'#�cI�����F�罴��$����C�k)������l�J�mq6�#g�3ч�jd��/w��{r��O0���I�;�����ޜ|�X���CV�\Js_b����ng�����q^�3����4�ޘ�y��Ѵ/��vH�H�x0&?l}����'�Z��&V��P�Eh��@��5[CDR��}�賹Q ���(n���� &�
pe3�[�&��1���*���{��l��G���
�ܶA�GU���R'�	QZ���oBtc�j|��Ԩ!۬<�h�sQ���j���"r"R�NWb�t"wgL�G	?���i�s� �/����PQ9��e0K*�I�Ni��G<8E��tƈ��6�w
Y��Z%�1������O����&����]�\磁�$�O�]؛���(��L�����>�i�\kFt���؆�"��ؑ���ճ��C���?B���ה5X��NO�nT���`���z�Fז�S#�������*_��Dؠr������M�#ri�a�fe����1���	�F|�uU��b��G���������_dN\��0,=�?��n�S�}�h�Yrc�;q�{�����u\1�+��A���럺��P��E����t�6i������f\+l��{�6N��_.���so-bյ*�\[id����bр��V��.sߺ1���"�[��q�W1�� }��N��}_C���C�P��?L)���L�F��|���|��U��5��P�*����\�@wn6���gm��ʴIT���#+ �t�,�T!4r1��T�`�1֜0ְP ,�����O�p�%J���-}���.OT
o�}�ru5O�	�4a����R1�my@��
J�c�z3�_�s�����B�ہ����0���QI��51(�7+�B���t�Td$y�⸎�!�Q�D���0O~���&3���BǦ�
�	o���d9l��veoT���/k�^�K"e�i�`L�귊�Z;�w�~^��_v-<"�KI��	x��55kv�壙U��(����BZ��QZ�~o}ӝ���I��Lx�	�/7ERJH«`	�FN1����^+��I��1�G�F:��㧎��w�;�7�ǊJ�TSNbL���/zY3�d;�>!:��5�#��2�Ǜ.?E�Z��ie�3
'ei�� ?B��Ǩ�j�z``�F��BE��58Y�{%��q�%��4���  �.�'�?R�ۊ��f�&�Dn{�E֯�:b�����R����A`��ӑv�Z3d�^	�(r#Ex�E_��0�M�^U��Ho:_�hM���"�9���I�i�#�b�ɰ��Q&�����%q�P�mk�m��x�W�� ����L�~RL�c:��DE��K�2`e迬ߓ,�=�c����Ʌ��Cv�x4��]��fP�7-@�.p�����4#@X�p�k��~5t�UQI4li��'�u�ř6x��a%��D;�.�>��~���T�q[���஍�i�F���l������܀Kk�"2a�8�L=I�}�#�ݯ�͓]baγRg���H�P�)�s�����#�-���	�U��/(>�;,����c�;p�̶��*�r5!M�c0�Gl�1Wg��A�
��	l4)lq!9��<ݨ��^7xt��e;�e@���U9�ry��|4�_���jJu�16�G����]Bu�u�0Q���믮���\k���i��9�W��%�eM���u,�[ʂ�șȰV@G�<��z��� �nW)ʢ�B���P�myK3����^Jt���,(W�9XdW��9
X��J8�7q�\~����˰l�O���_��o�j����������<6�D��)����E.Y��3�� ԎO���D\�ڄ0�j��!�f��X˞Oa��X���@cg�+��d$У;ьp�#{ �����4��r���A�˱�RTՒm�7/fZ���,e#ES�-݈��Rs$�Io�'X��V��D�|<^�U�<v�X�ʔ<�i��ؖ�/& �Th;���O.��0���t!���ͷ��c2"��'/ �^4vk,�`jj����tHW�g]Lx;��a7k�\������Ρ�	 �R��p~ �\��j�&��sb��tO@u�u!8ȦG�X�D�|�h���!�2P�����Y{�U=�`�h���M�yh��_������S*��z݉3K��]ƾ�����틺�����塚!�ۻy"韲�2������~��p�`ܱ�9y�?���#�i�qE�߭A44��Ɛ�"C��v���N�AA^."3�,��Ĥ�'���	yN�S�,�-���;X:�\ �u��5ԚS #x����{��ln�L��Y�������JQ�UZj�O�yJ��u�t�/�I�%
�n
"�a�"��T��GR)��yuL/��$7� 5��\bN�5��Ex�kPMQ�������N�����@����i���̘+򟘏#={?_
�vŝ�`rY޶��;� m)�}��]_w��90� Bp^��չƆ��M���v�G����ҟ�(��'��?�8��ڎ���	�)@������}���F�$4,|�)+�iLh|��)uR#���w6zv��jK)NX%�4��Q�� �79i���*3t6���EVC�������)l�}�c�awĔl:��O��:��t^��:,l�O3+rn�kↄۑ�L :ͤ��[��!RYG-h"�]�}�U�Ĳm�W�hr���٘"���������s\��l~l�yP$�j�:����g�N��a ��@j�"���.N�^��Q�k#�rgU���9J��>dKP�v��颛w��"� �n��C��sI��p���*40.W
�5�_D�Vg�e��}A(�q�
5�`\�d����)�,�hl�O���%K��]��_����6_���!q�~��+R�@0/��"i<y�u��r"�ȱg<��x�����jP��:�6n颇�/�Yf�~PG�A�i�%��X@JĚC�nJY�皲,y�z9Ͻ<&�?	1��N��mb-S0�a���}��!�u��[O�F�1��.�[���,P(MM)f�=�q�p���QI��G6�[v��> ��ܺ���J�IJF,�^�)hDdء��Wj��f(���am���9��n��2�(��ȿ-�ϵT�����P�§�*��&��=9W��r���/ eN��T�+�� ��n�N���F�7�9����9��怤Q����`kl���$@�l�`��6y5���A~�N�[�\�>���$�k���"����%�y�T�9Mv���ܭ���7�~�^�i��(����p�������n5�����(B�ӕ���QW���]TQ |�M�<:��M�c#��0ϫ>�O*Pf��[���<r$����Ի&"Hb!.���뵲��(̦�3���W��� G�b�&�j�va�N�~��-O�'�<E��r|:-V�9�i�����Tc�$S=(ص'^����"�]h��(!�ch�I(�V�*�3���2��Bo}�`Q�<����"hW���� x Fi�!��+�`CD��(��=�e�eo�q<!FG_��oS�J=\X�6��9ȏRg���Zz�G�����Qa	[���s�S�tӂ�q�/������r��t�ut�)�l%R��0�]q&D�n�\�w�*'�`��<?Y#�3��ӍHuj�����
���� ::��2�x��Ur��u�tRip�.a������M��S�,�d�5�_�U��#����zS��Tz5&�K��}A�D����I�v&cԬ��_$���jtq�S��v�vJ����;z5��Up�>(T:��G���0^w��Q~��5���'J]��|֟�Y�{{����'��D`°Zp.�R��v�#�D�P�����d����/������<t#�ח˗�h��bm�y�#���~����F] ԙM"�*�~�gC)cR���nNGX��!]��5�v.����ޮ�?�r"Y��۠{��~�h*�y�Mը+}0���	ڳ�kw��s���2��N0{�;R����Z�f�[ꃚ�7~��B1"Dt�|��M����=����:²����Ϛ�� ��x���
P�X�+,�����C�zVb��?���'�,�n�rZu��e����a꾴��R	��:�`%Ӱ^�P}J�?�����tM��ø\�3����S�cV堞�/��
�h]��aol���3�	�ڬ��{x�*S�g�3�^�3Z4��<��;�y��#�^g.+D��ΓmM��}Q�ɗ�&����PfH�O�p#��D���pXBR�>�����+���"�Y�$��f�]Y+��[�b^�g�ԣ��kۧ��`�|��c���� D?��8̹d�Ϊ�@ b��I���P��t>�R)[1L3L>p!/گ!���	['�K5ÉR��t�A�\=V<`C����1�6��O?7AIA�#3��C'���W( �����m�h�޹
C��른�r��R�{�i`���s򺢙�5L�z����푱4F�Ag�y�ü���NJ��+u�D7������:]�N�R�5<dD̈́�|���r�̣�9���hYڮ�[�cH<��b��NW���W���ry�0Y�`� �&j�r�I1�m8\ a�xM������>ӝ�~FG�P�������=�i��/��0NӚ�b�y�Ð76��F
�K��ؠfG!L%��p���S�����g��������O"��R) V �/�a&�e^0��wEɉ�A�fg�-�&����g?7���`+>���pR����ڨ2΍���F�u�r���@������K'�2��+��B&9�/��)4��6'�f��>?_#����|
�|�Ѳ_Z��~�X�����
��<�7:���Oݘ�3_l�򋟓�Vs���X"|0b�gu��+�g��o�-�*dܕ{�O|���}[ �͵������Ef���29���/Y����J2�p=���Q�Y��ho�ټ93S�Rd��^@'���-�5��B@s�O�T���{�|!���A��ag��b�v�V���>R���,�����Zy^�)�}�*�1�b�7�q�� �|m/LH^������s�i�@��Ԏ`�	\�g���  �鞏~�ܓЬ/�c�Rl���~'�.;%��5�dS�}�Gԏ��A�^��c*�&$W��I�Sm�	�	tUkB]�D��Su�",�k`�RAcw߱$�S�B�a�7�h��D����T�uN��-�Я�)Hz��.��9����F���YU�!6Sr���`�����C�RGd	��/�T<P��MJ�E��\ ������m�υm������VN�JJe�Gԁ� 0m��Ktd�v8�L�����<)ӓ��%;K�d�c����ip��ș/g2�%n��U���J�Y�	8�Ix��Wޒc$���ѝ�͚>Q��F3���?k�V*�&^b#�?�Ջ�N�2����5�mi� ED��˵��'%8��'i�t�έ}O5+�jg-6��J-l���w!'L�A�eVҲ*0�`v_8/�x	kV�Vp�u�҇Pm76~:�Hh8I��{ih��!Ҏ�ۣ��Nu�{!9+��He�͝�n�
Őɏb ���%,�hNzՔ����	]�wH.�D�{M=B���M��z��!�c����#+�����η�2i8� ݹ��~)�ێ�z$��֠�|%��9��T�u :)�X��GA�5e�󎄸&AK�R�f1�D��R`��ЩͿ��uWiM]L�d'}_��!.�X53��f䐹N|�j3T(����U���<hQ�����N'�;�$�����ɇ�I��+��������@h�'vɍTܦ����Ez���{����펉�tL���o��r����	������*?��R��B��2p��=R����2�
��E�r��ԋa�\�KMv���Q��VM_��� ��L�I�ᚇҗN�m|W�_�)���S�E�r�:�y�Z��^|_��Gʓ�T�6�x�!��l��60��ρ���S�x�V��b<7��`�"�I�y�O��!��<�țG�`�x�̔�����r�v�/42�]G6��sR�����H�W���b�	0qMV��X5 x�ܭ��_�˃m��2jQT)@<Yw���>y�������7��zp���L�6��U��q~^X)P�/��wCݙ�Tq���Q�e�U�S�)K.D�lvN���<��Y�}���_�;u���$�T+�_�޻�Zm��Ȉ�ȫ��G �|���s��R����z�=w�MP���<�U4�_�]����.�����8х�3
~���q�>�hZ{�ŸQ\����M��бcN9	L�߽ZK���׏�`��P�^�D�$r:�JJ�Wx�-7����ܔ�mq�lV;�Vh��J�7�
<�vc�� �z̓�s4�<�:�Z¼��5�L���P��b5��yh]��L��P�7H\;W�fA)�~�X���32v+���ħ���db��;��)�)����6>�'NE�������pw�f5[���nq��9Z��6)߿�;rB?��`�v|���\�Z��µ�,����Y�u��Yt��&�C�_�K%��ۦ��/�
�@�0G��S��@�m�.-N�6]��n�8�'6奛�qp+ݼ�?:ޞAL�e�~jh�ʠ��w���Āջ�C.�M�=/��5���]�.��[�ms�B���ozP�`,b�h���}�G�����~0�0�� �i���"�cs�{�8K�T�< �$N���bnb���P*4���q$�m���o�AСN��}��=������D�c2O�o�)�r,"���T7�%
R��pm1e��,�N��jQ̞�j.O�ܝ�)��Uk�"񖧡<��\���.�>�H�]�>����\zj9T���X}R��	<!O��Iר��F�����?�疟�eh�R���f���-4*_G�!Y�����!~|�D��ۓM�ȴI�5��~��x���{<����T��ɣ"�=�}-C��E\��g@%`�~���؟���M�X�Z�D�F����x�JVN��� ��5w�|�yt�SH� �Ā6���Ɨ����f^s:2� ���'��zX��u˪H���V�C��2U��o�Զ��'�=��2�%�_�Ї�+�����$��DiEƟW$f|�>�7I�G��\}�%�xQ�������Ǩ
�[�R�1��o��&`��^"]%0͠zy�mD<sD�����p���9�ڥz��D��p���ݭ���c;�G�9VW��dP8&�+�l�W���?f]�ȔB�E<��<3�y�,�h��+<��rA�d��D��\�W��<C�����T�W�z���m�%]<��J�H��w�+����5m]��~	��f�t4�Җ�SWX_��^���9�!�����ۈ�I���,��t��x;��DL��G7:����/:"z[G�#����i��SC^_O�����/'[�m��@E�AZ"����z@S�����I��9�<����̉!�=��|�anJ݂ͤ+@���lIyz>Y��'}�#�*|�S��kO~9(�&�E����u^��q�E�_�.<N
h�03J\�����'	U�=���w��:Ќ���
NN*�[��E���rX�\�L��1c���
���� A	f�w� �ՊH��y�@�����K��=�����X��}�
s��g�^#�R9ju� d|j�k�`Ĭ������n��&ĵ �rF!�Ă'�>_��\��z������T.�q���V8�:�~%nB9V���h��FH�5�g8�5�(#��V*NC~�IQ��k�8Y�>}~C�n��3m��
�^0�QL���q�D')4	>�X����x�
=8�d���bT7���l��Շk�*��]	�<�P�3�z��&H���=7=G�������=�	㫮,�����k|s XL�i=ᮁz�|hu���'�<��B5��V��$�r�8���[ޔ�(�߽�*�}ۓ�B���nodڞ��&��WE�g.��O~M���� SSlz�W�h���J�,2��S��Q<��؀r�O�C���;��{������y�ْ�����Q����Qd8:D�Z��Wn�� 3am�C��j+���6��r��&U��')^0g�)�@�-09=N#���WS�s�SH�l-����R�1�g#f�&�>x�{�ǫ]�w��a���kl����C�g���T0�I��,D<�N°���5/"��?x�Ac3NȓM�`�|(�,��[ޟ��++|k}
w_�8x�зՋ���Oq�̛QpC��h9�y}DS�4�}��;�� y�)q:�?w���D��xUi���%c�A���B�5`3�v�sD�h�~X��"�j��D6.f�v�p�"h��km�[��<IsY���0�ڦ��`��Y`�l�\)\}���sM9��]sK�+�.�w���)3�t\����K������naz
F�K� ���&{��4=As�m1R�l��{y7%�j"���3d�.��Q��n���e�<����Y�~408��:�^)3�=�uX%��<�>�g��Y����u����w:Y�S�
��K�ǉ�uaN�/XǕ=F~�v��͏J⊞V��A���V�����d*�p��w�sJ���~���Ü�!��X$}�K):?�/��jV(���))˽<<�+��;��R����x��6Q$��&U�b�<Ԙ��6����2HE�c�Bᥫڈ��1��v&�������y=���b�8[�@u����u�j��֥��β���M�R1Dno��b6|%�0L�����}�J犏ʄP�\_��dA,?����JT Ų�y�(p�BJUȚ�'�ۆX����}M-����U���>5CB�_�����߉�3��z�d/Ψ����\��r�۾0@���	�+F�=@��q[��^�m�W��"��#%���r�T�SHLM�S�G�Ͼ~$�j���4�i�;'�;$׾}�$�ߑ�]bB�.-�t��̧�fk���rM�z�h�>_��[RQ�
�Wͮmok'pC���m���b�7/�	�*�pAcP-��:����UH��f�~�5�$��3V�T�B,� �3���9�$h09l��~@��fw��T��ޑk0����5����{�՗9h��L�����f���'�Nk�Qp���]/U��?q�p%L��3�0�ڈ_���D�=�ٸ��D��aH�v�3�ůPJ��V����
Ra.��u��lT��������Yy�ئA�zwy�Ϣ�Z%E5
�kT�ы���a�x�8W�;'����/P���m��h��P�G��MO���#0���9y���񤍼��|%���T��jy�g�c9��d<�e�pn�.(���1��CF��mW��7�v�ۤ�T�E0"V���"%���.z��!�F�r�,���������튶�Ȍ9	vH���q�vq���:�����$�M pt���x?ܕ��(3H�oU��ߴ�:(ɺ�'Z�tQب\Q�%�۠G���3?{����\Ov�!��<��/4B�'OI�!s�V\�����{}��JT�?-; &�] �}'Ն�a)�����ܵ��)�#�f�Us`����&���e����4�.�8�yܛn�T�rT�o�u��h�����R�D�R�"�;��۷s��Ȼ�=���������O3�S}�c��-�J��O��m=� w�/ �A��:kW큝M$�Œ�3{�QK�,�L��,{p�(Y�d��>^��ꎨ��5b�j���Im��!']�ՅM+�+Xu�
�~~���z:>�����I\��$��zE��E,�Q�!h�h��A�DC�J�~�w�w��6;�vޕ�^�P���d��>l�_}f#���Y��d y�]�:9�|`!�wE�C�1r䣺VO��`m��i�9�gGh�{��D}s� @����Q��tQ�����^���Y�:�
���r��in�X�	Q�����^�,��V_ѕ3��F`�I�P�b��ȹ��(p��X����k�:��
�%z�O��c�}[ĮC�d����)dx��b��ZS�+�6 \��ؽ��iX��d�!�`Q^��F��_9�L�9%��#ݒ��#^�J�x� Җh��ϙ��y]����JfS�h�A�:�&�A$�W|�s+�wx����k�N���p�����P{��IB���CJD:X�voU��AH
���y؎�
H�e"����&\���L�H��j�$��[���B���C@�缰[�c��[L��scXl{�
@�X���L�\~�݁:���bd+ku�ғؽo���R�����/|�k��ۡ�����������Z���g���IU���6�H��� �@t���^p���̥H�{"�{�
�� q���&��	>�<vw, ��qt�[���[I4�]M�UQ~(��=����nt+}�����Lؠ�7"��	�V��@�Ks�+��,���m}�>�;������9�9u���զ���̮�A�Q�Ě�#���9i�>