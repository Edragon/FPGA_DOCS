library verilog;
use verilog.vl_types.all;
entity altqpram is
    generic(
        operation_mode  : string  := "QUAD_PORT";
        width_write_a   : integer := 1;
        widthad_write_a : integer := 1;
        numwords_write_a: integer := 0;
        indata_reg_a    : string  := "INCLOCK_A";
        indata_aclr_a   : string  := "INACLR_A";
        wrcontrol_wraddress_reg_a: string  := "INCLOCK_A";
        wrcontrol_aclr_a: string  := "INACLR_A";
        wraddress_aclr_a: string  := "INACLR_A";
        width_write_b   : integer := 1;
        widthad_write_b : integer := 1;
        numwords_write_b: integer := 0;
        indata_reg_b    : string  := "INCLOCK_B";
        indata_aclr_b   : string  := "INACLR_B";
        wrcontrol_wraddress_reg_b: string  := "INCLOCK_B";
        wrcontrol_aclr_b: string  := "INACLR_B";
        wraddress_aclr_b: string  := "INACLR_B";
        width_read_a    : integer := 1;
        widthad_read_a  : integer := 1;
        numwords_read_a : integer := 0;
        rdcontrol_reg_a : string  := "OUTCLOCK_A";
        rdcontrol_aclr_a: string  := "OUTACLR_A";
        rdaddress_reg_a : string  := "OUTCLOCK_A";
        rdaddress_aclr_a: string  := "OUTACLR_A";
        outdata_reg_a   : string  := "UNREGISTERED";
        outdata_aclr_a  : string  := "OUTACLR_A";
        width_read_b    : integer := 1;
        widthad_read_b  : integer := 1;
        numwords_read_b : integer := 0;
        rdcontrol_reg_b : string  := "OUTCLOCK_B";
        rdcontrol_aclr_b: string  := "OUTACLR_B";
        rdaddress_reg_b : string  := "OUTCLOCK_B";
        rdaddress_aclr_b: string  := "OUTACLR_B";
        outdata_reg_b   : string  := "UNREGISTERED";
        outdata_aclr_b  : string  := "OUTACLR_B";
        init_file       : string  := "UNUSED";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altqpram"
    );
    port(
        wren_a          : in     vl_logic;
        wren_b          : in     vl_logic;
        data_a          : in     vl_logic_vector;
        data_b          : in     vl_logic_vector;
        wraddress_a     : in     vl_logic_vector;
        wraddress_b     : in     vl_logic_vector;
        inclock_a       : in     vl_logic;
        inclock_b       : in     vl_logic;
        inclocken_a     : in     vl_logic;
        inclocken_b     : in     vl_logic;
        rden_a          : in     vl_logic;
        rden_b          : in     vl_logic;
        rdaddress_a     : in     vl_logic_vector;
        rdaddress_b     : in     vl_logic_vector;
        outclock_a      : in     vl_logic;
        outclock_b      : in     vl_logic;
        outclocken_a    : in     vl_logic;
        outclocken_b    : in     vl_logic;
        inaclr_a        : in     vl_logic;
        inaclr_b        : in     vl_logic;
        outaclr_a       : in     vl_logic;
        outaclr_b       : in     vl_logic;
        q_a             : out    vl_logic_vector;
        q_b             : out    vl_logic_vector
    );
end altqpram;
