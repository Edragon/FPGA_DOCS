��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n���O� ը�fN�ݏ ?b��[_�=0hK�v�Br|n��vW]�pz~e�e���O�Qsv�g
�i��H�@�yޒ��g��A�mxp���I�Qt��Fm�ݾ��CˁWfaΚ���>*���xwt4��}�����z�Ê��̕H���Bn�嘞�%��qF�FJ�I	��p�v���q��Ѣw�Y@���:U��C12�"�J}�c�o����L]��ALpWpv��ʸ�-�r.λ��-��hoL�!��]�a������#1�'f�E$�����X �2��^E��&��,�FJ�tC�F�_�@��ݲ�{��ٚ��ҵ�s��<{6lS����)���qH)!zf��U��ޤ�N��&�-b�D�NᚆTvT�2h1�m׍@�q;Hߺ�`�gU���GB湄<޸JU/�O׃���߳]�3 *}�Bj��mx9�n4����b(�Y5
]����"����!o�_�a����R1э��dvD)	W�f&�-��g��ծX�.�z�b�SmT	ɫ;�o�\�L�(��	�s��;O��U �	G�#�ըz�~�Ga#wĘ�Ϫ{>�xfe��u�VP�&dje쪘�T�����
�n�Ѫ*p���3�.3����̳��y�����-�F�{�%���7�+l�0�0����~o�k98R:.��|��m,��9�K;ãp�j^!/�~<۬�x����y�!I��*�q
c�m4]�+݄�i�qK��8�� �Vޑ�;�D����8����b�H�I���g-�jo\��j��Ղ�Ƭ �-�n�lLn���\����P� �ǃ�]�%���5��@��=CX꼋Ģ),��9���1�B���=���?P7��C�ls�7����8�7=kFR�M�($uӨ-:��}�R¸ױ�0=��\>�\�ܢ�9yq���s���6�x���5/G��K.U��D����1׽7p]O�@��Ș����:'���ϛ6U�|:[�%���T��D�·�a���jR�}h�ג�q$�ԕ�&W�X�o�~R�8� uj�ʵ����5dU%0X��7�n�"S���#�P���$"i�
.�w.?t	V�Jn��]C����vU�+!�4�/�"&6���*vh�]A+�_FG��Σ����n=��=�{�'�ަ��e�o�k�a�t��������n)��z��7���
��7>�	���'��;))�ٓѾ��҉��E��	J�;��d����3I_|V��lT�1:�"I��!uKx�Tp�_ے��p�n_L!4��uW�J�RA'�y�x���ŵ�$h*��?��hJ����hAA)U���Ժ]
J�b_���Ll2�@��ubEE�6^S����m���}1+��;�3/pg�e�mWQ��yW�"���VL	�d�l��tA䋶O��J�Фv2�c�e��M0�8���� %���U�_r@u��o�;?tZU����kX�S�	�(xS��oЊo&��p8>����}9q�*��?.�b���B�Y���?�ȅg����f��-�'\`HB@���_�����a�7�F��Jw/�bcM%=�T�"Sz�L�5�IpJ]׎F� J��YchQ;�
��|M؅�^!LW����k��R˹sH�	?2Ñc��ZgW���-e2�и%���^fG�e�(M��e����G\e�c�R���Ӳ��K87���r�����"�DlhΔD�9����N�m`sO�}��B�����;Ko�N���L��a53+��p{��n�Gy�tm2ՊCh�Wx[B���,p�s��D�զ��=���p��\Ԛ�̈#�d�v���qf�E��[G���d���)�dM�g��uI�gnX?�m������2!�(n79=���f�� ��:��V�Z���f��Q=���J�ZV��,,�I�t���`�cɧ��t�;1e���������*�Zs�>K(� ������S]VQ��D���٘�ݣ�gI4�c����am��T�Y&^u>%���_'��&�h�JaK��L�ju��1�d�?�����E��ﵺ~�
	� ���m�(���GU�l���n��ױ���{�w�O��k���d�31Ѡ��H2��`HL ��L���)��vC	s��-^V��9ǹ�2cu�׶���x�l
2�^��>oȖC��ё0#�k�uV�� xwQK�F.~Yh_��4�q�*;h����W<N�r�v�yc��:Qu�朓��0�"�Q�EO���>��>�b5��v��'�(,JoxWE�16���˟�\?�k��&M�w#\�j�]H�|Wlh٫]x޾r$��ڡ���8\����@q�hO��~1L��Y��X �t�+�3j�i,����8|ƴ�y�؂��
E{L̐�u{�FMC����}}c�Kw,�<ͽ�^��3e|:�ZJx��h�"hjE���\� �?p������NG-I�oRg7��-*.6�:\̃Y������B�u�΅9@skQ�<� ��1|w����oEN������dۇ��>|�Q��7 \d�����&�j�Xێ�� �/�$�:�VZH�\s�%�Ӂ�*���`~bQ��<�f�]��,�e�6vO�����"O��-���!�I��t�7n�"S�~!��M��b˹^W�;���K<����&9���q���z�a��y�2��(Y���lo�x�UT[Ŏh���@&g�o�P�@����N�;���~�=�f�x�8� ��f�T���d/kUX�jN�5T��[ӟ�v�+�"d���{�?22�)�-��~�u7 �(�5��i����*��-�p�����J�X�B_��K��NO�B���AQ�=���si3<�R^v[|��>�7�:�OU�<jt�� ��M0����쭩z\H	Y{9�@s�\�j#"&�~<\1�0�j+�OK�N�jn���4�r8��j�A�w��$궏����A�����5ݧ��3,c�&%bi2R��6T��6e�N@���붛��ɏ����GK�*4#^�r�P�^̩���-�Q�%z�L�Wq���d	����[�>h���i��m֔1���m����ǣ���S3�/�	&�WA	FW� �T�Sn�Ӕ=jK-�v�*
潠�ʸ��˓ƨ�� t���\�ml�*��b�$�1��7��]��p��m%�*L�(2 ��{W��������o��چ���ǟ�MGo,^v�B��?lJ:���;�\{�s��� ����5<�q�ĵ����ߍd /�W��'V'e�����2����XL�V5��qW���1D*��=�k���\<}ާ�W��	�h�-�-O���j/�Z��!5�D�
��B���P�Z4e�Ĝ���`�kh�37=�9�ua}��+�~e�@�H"��b	`|��#��π,�r�ܧ��lH-��e�s�vT�F�������$9T�����;�#���}<֩K�@r#ͧ�eش���Z�Ь��Р��c���ՅV��BW�ܠg�QI�ŧ��S�,�£(��J����=��b�w��hX>P)[@�؜����vH�j�?�$tmai<֠Օ	�I\:��� ��-�d�J��8�(Or���X@�!4Ӎf���Rb���	E=�Tl��f���.�]Jw�������������Pn|��x�G�YGKf��OQq�nk5��ßXV�b4��2%NL�x�y��ϗ�J~���Sן�E��8zir�K/+"�D��`X�H�l����_*��1��]�@��l���AD�ب��]L��G��q����r��3[��yZ��O
~��:���y�d�i�|#��<�ݩ����{3� ��I�a��n�yz����u�����s�T�Tskf�����3��e�0�yJ�^4�(?�XƧ�_�Bԣ�#�BAF�H�G�!���
��R�A�<��dW���$X�=���q��S*Hƍ晐L/�>_�!0��+��	jh>�>���z�{��C��~�Uw<輮+���ݪ%�f�6D曫��rc��~��h$)�0������k�!��u�T'�D�wE#WN�F�S�V쬚����)�,���;�l����E��,���װ�QTnQHb�$x����F�W�;@���	e}�}���H��L��Wϊ����� �����E�k0���fl��OB~�y���s���������d���շ2�v��`��!�˟�:+���j[u�i�ے���J�����BC�1�f"��!��B��9����uۋ���r۽6�8���4�˙DK�O���9h�����8��1Ra�O���|�4\�g�n�i�G8�z@�<�BE�/^ ��g|Z?�;��,�[SK�}ς��ԭ���@b(��_�<`μ_!?�	�%��̑�7ޮ���N�r�!�v�&�X�{�i'�\sN��_l��Y:L^ ����~ ��m >QSo���x�'�,t
�(����8������l����Hq���� �w�8-�Z[i����$���6��H:��:���0v�A����O� a1�x*��TW��
"3�\۵���uK�c�)Ǻ�1��I�!T+Ig3����Oy�o�螙���¾���� ����X%��c��?7���v8�TmH�(� �=��H�`�]���eL~�|s�2���D��(D^܇=#����m7�sQ Y
o�ShZrA����"�}���-
T�����wgн���٪Qb�gc��v@�����/����h%�
)ߥ��{��Qb���& �lJ<�(���w��q�誤�Ѵ����V����j��s�6���6Kq�h� `э������*n&z���BZ,g)�t�=<-�5�/���iH����vqK�:�CO��:5���Ѓ�Qs��.�-�6���ݙÿE�?�^��x�=���哦�/��!���D��1�2*e���z. ��9q~���@��OK��{����u� J4ȃ��+��":2�"ځ$2l���GW����Ew��縨Ú��c��~�I��������}l,�� �!���VHu�׸��_����Q��Gk�X	��X�*��oE|���َ��!V"���Ϙɐ$��&8Q�M��;�&��f��9#�f�[<�$=��� 0m0f���ߩ�R�ūɵ�+��+��E�W߾� 2��C�h#�8S��1�0�S�]N�wr��PI��\6e�tƹE�f��Ӭ!��D���ol���W�l�Ф�\�Qz�d�*�e[N鮲 �ӣ��zq��䤂��(1�ު:v*���������!|�C��s�IDll����M	*s'"��g�IZ1h�ן\�?	��x��v��N�I1�΋�,0B���ؠ��g���Z��� B�A?6���0/%�7�9�ʰIK��AhC`%}\��ց0� m��Q��R�/���$��ܖ�3�p�~pD'������N	���T&/��bd�7|�R��g��aMT��j��3{	���k%e�(m��,Ȁ�R�<���������[�P�k�;.�v�=�߄U
X`*�j�1�3�5�0�)ap�W	�V���iZr��,\jJe�&3���\�M�Z0_��m�7D�g����uO����w7�/�^�~���)e/��o��[��q%��aTZ՛����"�e.@���aH�t�w1�b{��ԕ?��J�r��%�N��E%�LL���G��ypb(6V�-ܷ�c���i����a벱���QS���J�Z�i��Z� }"B�~
)LS�X�?����J������=��t�Z�_�b�N�M���{��&H�*��妿8�����
/�E��1�'�a���-���}.dxs�0]S��7N��y�����(��EDx蛢��ca����+#_}i��y�h����K�2�n���o��lH���'77��ɜ�s
<�]�Ϟ��B�i�Lkz��M�0Q�0j7  n�F�h�O����Є��j��빗�<�����?+.g����5Mp5Ƀ�$�2y��뀟��,&��g�zN���U*�h5�p�X�m�� ��ֿ�ȯG@ʽ��=�&�Q2f�*�{J������ �>�T��;K�U�%�]�t!B�4R �cB"Xr��ҍ��]kp\;���i�$�a�.�G�����넇.��(��5�\RB\ ש.�y����{��!4�7&���w�����Z��n�� �)�|7Rx��f��靻�ڎ���b�"��� �̉��X�"�\�,2�wM��{U�P������Y~`1�_��D�3����}E`��Cs�RQ��y(�J�l��Y`��O�1�n��9�3�P�ce(}u����?�_�VdN;�gg�ll,��[:w�gŀ+?�X~`Z�$����*!^������Z'`���C�G���v�\Fv.;x�YDp2�`�}�z��j4)�̗�z�_�<N�"W|��1V���f�\�8r�Ż�L`ګ���Q8�����V���ĭ��b؁T`8���ʒׯSH��~L��ؒ��!���n�t��l-yy۩�E �|xnZ���G+���q���b�֞m���,֯G8�,K�a�0�,$�9v�� ]�}�#����{�x������u>j�zٍ!�p�к�Lʉ�,�W�X�n�p�=���D�'t�"�Ķ�p�1�v��J�6�p�X��Є��d��݋˳a�_X����c��]�l���Բ���H���U��`(���:T:��-��%�=���&Ej'n�
��?e[�'7l��S6����¥�X�,"���4�&{*]>�=M_ huUu���^E�xL�/����e�ܥ���������p��#(���j�o�2Կ��C��lG�d�1U��M Y�� L,�r��T�c*��D�[���SZ�S�ŝ4�X�3�~ʧJ�K�����	���$�E���(���*l��)�F̅o��� p����C�Ν�����O�,���Ӊ*Q���2���(�SYS��#�����Y����x�J9�Mx�}+��;.�d��M���W����*�\<u�G;�Pt��~�Ӎ�Z�;�eEx~���f_�DE�� ����By��RSJ��ջ_�h�a��� �=���6�G��B�Չ,��G�^1�ƫ��Z	7��G�S�����%ָba�%������Vg��iz��1�i~�9�N�ڦ(��5��(�r��0Y@�y���̦nY�}iMq~O��Tm1vhOD��t�!��
@p핪� �M��������ƃ�SHb��cat1�<�����:�Z7�L|r���}�H��E�yH,��Eb
�Y@xOm�f#����u���؉~�q��%N�5��1ǿ�0X�x�b<Xp�xd��m/�����f�s�[��~�c�5^�F16�C�^D���,O�A1͐�}?��#�v�5����oD��0 H���uLs�m2��K�Z��Y;�BP�\CQ��뿢�<ߟ@ݲ�9���'<jŏ�>8�RpȠ�������ӧ��Z�+�ݜ���A��n�'�� c(� �}��\��:1��a֨j;2�=y�z��p{
���X���ګ���(f����Rʠ��͕��t����7��<=�%_s���N�,7�5!}�
(���\:{�Sk0T�E]��l6��*�������>q`2@}yV�C�Lk��)�У��ץ48h��	���`P�D�Q��4xB��	�\r!ΐ���ꁨO��Xn$���+ޟ?�d4l"�u15�zy�=y��8�̤��E�٫�@����g�
�P�2ga�YQ43����
�{@ץ���^;R���o��J��k�9H�D�ƻ����0J1������'�i�4��2��t	V��
г���sk9Ҷ�]B�;���!o����i}%o��:
�H��>Qw�0�nJN�ז��8�D8��:�{�c��F��}:#݇�͈��t�N�z^��G��>�����N���y#���Ո����7�R x��B ���!@�KD�I�sq�E��a�t�:�K��O��A$�װ6�eE} e�Wu y��if�NIx�uU�oX�{5��qj"ܔ���E`�-e2�q<��*����?�G���G�z��dD�t{F�'j<�V�:���|�}{\�h}����\�{���4�!ʸ$žx��G��{>�z�{9\�����O�;���Pҩ2d�I,R�
�C�,Uw��ߋ��?�w�x�A����|0ގ&���i�	�'W�ĈQ�Q� �h�0��v��b����%�N����,���Ɍ�����%�O�IVFf�)J�B��~ }iҼu)�vV̈���Q������-p�6��dj#�-O��ʬ���r�m@��%~�ʸ��!]�}�wqaYR@�²Q'�d�]RKY3���E=���\v���r�8�݉r&�B�T�;�סw��U���*��+܇���A*�!��O��٣��:}dP�{���;m�3ʋ��@���#KD~M�H��jt�p^�=�A.�ݝ�>����|��/�����d��zߚɠEscS�������vl��#�\�L��i��\Qyx֞	���  �
�D�:Q{��4�lҫD�����3;�,v�e��bK
�L�XJ�4�۹3�S���cK��Xā��I��t0�b�䔎s��

O4���#;7Gӗ�y������o�%���o8�T�<��q�.[�Q���խ9��F	j
2=FX�d�Mk�&l�ޱ�T	�!��ХT�6�H�l���+�]R��0��Edm��xA+kv��;#�Ru��#E� �,��G�!;E,�ޒă���Q����>;�Zk&{����j�f������S�y��*���qԧ��N(��#|FQ�T"�����I�UgU����� ,�]�4?�F����*��I6��x��k�nKPҀv�`䆻Vс ��W�c�#��\���UyB�"�y\�2�?L��."����[�٧��V'�	��!+C,j�[Ѕ�Ba��;ǖ������?ü�N�UE��
ɼ��,��@	�UX�kE��&��3�-Kj��X����S����w����l�w�h������:�_���������I �=>$��c��*�c������*X�O�A���81��G�P��wA���_w�3`8m?,�� l/��YA���b�x��VI����]�9qy����}�r>�^�����yL��y8��<8�K��V�g�����,����X�)�r�f�-����	�NF4�&�g�r�*��#�X#�y�g�1J�
�E����_�q�2g�|#��C�R�w"��@�Bt0QՌk�p�g�wƦd���FW[��h;�I�����$x�2>n�|1����Ga
A����$hx/ެu���j�W�t�iι��i��gK���_#��%�ݔ�W��yg3a�`A����G����Vk�ʺl�(z�_r��k�~�7C,2j���Z#�9+��*V��m�e�b,o�����U��~�����g�nH,}ki���o�7
q9���*bRmo|�C$�Ma��o�u�d���o�Yp���%�pX����c1����$q-dF������u!F�#��߽I(��#�}�������G�� Y���Al�4NE�5��6d\ˏ��S��xT�n������b�c}?�i��.hp��)-j�Vcw�3̓��Z��a���f._%���`�B�2$L�����:�fZ��l��߈w�+�T����7�ư�2��6-������X�����9� L�@����n����'�l�
"�s����ݬA�bO��0��*+i*U�(�h3<!4$�f�Ɍ�m�ς��WC6�+rN��v�q�B���Bf�@�x&,�2�6"���}un2Oh=)�^��T�fǽ����pFb�Ƃ#_Fk6E�Y�f������{����L��k]��h��1j��iV�]�X�r��_��^�,H8J)�FÀ^�OE�҅��կ�������:�,��p��9a���)b��x�D[M�de���ˋʉ��?�%d�BR?�g�����|��8��iÂ'�.K�=�%��U˔�J��=���CYZ1t+�n7	}�qL�*�	A� 9-�d$c�<V���i_'�l��(�vfB�P����PJ% 4�:��W=D9=N�<��w���ͷ����	�I�?��(p�
�6J�e����ݷ� P�q3�������	{#�$��і�\"��E^F ��.x�\�!tHb��۬�B�/��Kd�M�p=r"����RT�w-$�SuW�3+&�QY J�"ӭ��^%v�)ip��\Y�֐`�W]��7�����L]	���iC��[�g�$D`.���3�jV���G����*#�w��.U|�����E�,ƣ���a�+����UJ�4��bn��{���Y��`�s�� :lg�G����A�H����yC5_�S���|����1��IOv�m��F��=~{�3t�5A���,w~5;���=Zk�Xs���h�1*nj�.���845�f�O|��]M�"gLjD�l��y@-�8Bg1%�w��^���Xs�tё����Ƅf�=�6U��\O9�ǥS��{�%�$6(KcfT�w��u1���&km(8!@r���\QbX�",f_���|0���E�j(s��P���7���B�n�$yk��J]��/v�î)��k�@Z���y��:���z8x�a��盺7G�ɸ�B��`�(xd�2ďv?8n���h����c]��J����s�ަ�P��9<�&~=i<)�"�-�(?�"t�c��pa�Q�b�)����ܧJ�'}Ů^����۵\�6�9V����PZO� 6/6��|.6���Ii�X�r��8p'[uKL�h4�/R,�w�T&/�~���*|m�K.�V�'4���[�8ݵ+$��cM���{�L��J�Y�Jh���0H��i�`'��?v��O��]0�o���Ʀ
ڝ�ޅZOT��v�t\6ί=10��7�	>s��~���h�p���x�~�J�Cx�.U�xf��y��T��k�.��l+.��K��O�] j�\a�IB��@���ĂFS�[�CY��M&���a�fsql���7��a�%�Ǟ��[�VtS��O��b >�X��Q�J�sw;�a��O���C�Jy��|-w8�TH㾹O�n����F�_�6<(;���zcyk�^t��+�o�R���֏Rq�I�EX9�qc�iɃ(S�)�m�%xc�h_m|��lF����b�qb-���J:��2Vy�Z�M�����?��%/��RT����
��ިDsp|�y!� �φ�u�z_� ��*��)uU�O&������%f��0v��e;�k��JVq�U*�_+3��}`��"�!����C��Ƹ �]36�>
t��N��|�����[�������>\y1��*	�r��{�k''QRw5jt����6����LOs*Joit؀�C��>�:-(F�*�wWȜ�Lx�s.)���,��?�#��-�u44�3MR	)^�9�D�M�{�L�0��� ]�D�@���O�`�b�q?�뤓g�f[���������O���8��5`:�;�p)Y�;�ϻ���@��^\~����z�)��y��j����z�d�5��}������
7(�`ӂM��c}�^��D�l~�=)�S���(��e��G�]5����$�(���aM�7�L#MHC�>�����s�����ڣO��u���Zk�걞J�k��+��Yr�o\R!ٗ)� [�#N�ø �$��l���&�l�M>�d�3��z���|��j�M�k��7�'|_��	����e4�R�O��>?��uA�=���=a�����61� /�D|����߆}$f��Nx�^�~=2�������ƶ�:H��Z�?L
����*�Jd�(L�y�m�p�oJb��U긖�#�I��~"#>���|���G����4c�9�R(^���u���ޗ�-ŚENv�1�5�U5�sFl}�����(�t��x8[��=>s��a�MD	���Dw8
�����(�\ֽ~Xo��Rz���� �!i�!'h�<Ś`�bT�v�2�0�ܲ�B�^H�y��I��b:�����������8�� os�J���sPuw�)g��%VP�!<��u�o8��Q��#^��Lu�1�f}�L�!���GFdM-�ۊ�k�ǚ����Sجl�*O�y���2s����Kt�K.;I樖�*[��ћO�v�K쓁vq=���M9xȋ2V�)�H���|z�^�[cra/��aS����U��6	��P�R�^������x��h�O%`�Te���ʼ������U�Jժ��mo8�`ti%��#z��%>��Y���܈ʆ�"������Z��'�=]A�E�t��Vج[��hra�j�GcԔѰ��)�q�j�@��*0w��!}���ֽM�� 1u;,G[��^[��"��yqPV
I�qE��4��gV�����Y0����T�}��T7��&18KM����>�<��>�3�*hU�򖰻}����P��_7�kC�vNo`��:d�>�=W	�o�2�O@�+�2���v)��.]����8W��NX4ف<������5����Z�$)��/�%�	��}�G��e�43%�\�v���e��-i����}�g���G����@9�7uԿT]��F�c���g�E�ܰ�8G�1��$����Hf�p�tN�DB�}7�XzkyqT?A����H��-�����+2�|+���'��T�5�����i|�,[AU�^Sl��3��g�:��k.�\YdG�VBg%=��,����Z�Ȣ��E�B�Nc�啾Qw�r�pO�3�U�̿x�pQ��J�hE�h`I\N����nZL����� �(Gc)��kھ<��T�\E��qe�$�]y-�:��r_��߅S;Z�%k�0�G��[,�����a�Q\gia������+��x�A��<c��JW���c
�ؘNI� n�)x��r��:�#�ɥu=�
�,�q�*92���ىxz��m��	l�=�#��h��ܑI�d�9��Ƅ��w��ߦ'�yH%DA Y��q}���u�=����0�w���e=Qc��x�"�(��PPA�2n�Y��d��q!'M"�Ψ¸7&���=)���%#��.!Ը�B�"��{7	.����_�&r���Z�*�� �[0:Sc�p�q�^�\L�@��:�t(�(q��}־.
\�0,�qW�q>@����Vv��źH		e�]k�Z��b0Q?�������dEx�=�k�.)ɶ��hA��j�H�Nk'�x ;����e���g� _q�lք���*�ͻa�w����oڱ��z��7mוB�������I��`����u�p"�g�E���e�`��î��}����o"J�]�ˤq����J����;E$*���mcʅ�"�C�.-t�m���0���&�j�I[MY�N�ȱ�Ŗj.։�Ƃ0Z����o>
�k�R��v��J��ǭb)p@jP���H�(0M�l2�����+D��
��%���!T��'�RY��)������'��m]p���M��"��;$~ ��*�D��(o����G��:��&�ˉ���B窱�������9�ә�]pF�?�<�B��+�Q{�ާ�H�����~D[;�2[ͧ�Q���E�X;)��s\�]�ݼx�4Y��K�9��x�
�m�:ґ�K�rd�y
m�L[�/
�[]�S��t��}����ɤd�R6.m4�W����'Ì��y�o;�A0.ߐ��p-��pgI�����@a��K���a*֗�HJ�+�I>�L�a���
��W`f��E��Sάu�
`��LE�l)H3
cM=��d�2�����)Z�H�Tiɉ@!�a�~D�C���;E�-ni	�́�ui�E���<��	cW��}�o�%p�_L�Y����aP��ݺ_F?<嶢Q�<*@%{f"Ud�7Б^n�J�.������p�"��lg߇M�On�?�"P&�J0Q�O��'b,�Y�SՄA٪�|�%E�)�\�Tw�Q^odݰb�h���Md�e��9��-��A�c$�9��a
'�S�{k?�+S�x�A�w�ֿ���%���R�+�9ZZwd*��1�#���x!]��Ƨ��e=3��3��.�P���V_��l:�8��OL��
c柉�Ga���$mt��j�j,/��4[/��?Oj�p	a�����~[�� ��5��R�
�D5�#qf�L����<G�wʷr�(�Dc�5�_tq���ţ��II{�c����m"0j���7!����w	t9?N;#�j*nM�?B�g�\��li�?y�D�/��%ԧW �(kA�Y��J�
�Ьi
���s��S%��jt�� �������uᷬ�	<���׸΂�xP{��H����4ヮ
28��ȹ���eG�u�O�|%Fri=�MeL��#�#{��"���&ӣ'qW�	9*��S�|�'��MG��AE��A맅�� ��F�@):����YTA��~6����	41Sވ5 �f��%�KzUڋ�Nd�by��,����<��$��\�d��W�k�f�������q������:i���P��mף���D�q?PbK��xb���*���qH�CE4����
2��)�Mv�^�7A�p[�=���rU*�gT�y-��޶����G���m�m+�/W!��x��!��]������ևG'���L����s���ntu'���IG���{`�S���Gu���2�7�q'�� �K���9����C��j��(O:E���N��={�`��r�� &�����,���CX��~$ZT�$�Ͱ1�7��x��LVzӆ�/��+�GKc)w2�ߕ�FHYJr�t��}
�T�$�)*\p�)&#1X;�n�G�&b�Fb�.�JM�@�'}5�O���Äk$M�^�e�a�_��||'�$��!�R�;g�[�(�����K¥�m�~3���/g�PV�\�Fa:_�&րtW_w����KLV��l'�bEz�s[ �����ƅ�:�@����q���I�تHD�����R�R��Pp��iݭG��;��du����O�0��**XRg�x�P��:��C��tKaH�a�Գ�؆7h�S����]�=�>�	��wr�b��rH�kj'��S��'a6B����z�Ʌ����K^��k�Z��b�vk��7��)�J#ɚN��O��6CV
�Y�Yf�su��ug��19V�������O�|k���ִ�`�(�I�dٱ؇��j� ��E��|�Y�"���]���h_��nr�Wm�3�)�V>B�;L	��ĉb�D�����0��gnZ��6c����w!�]eI9L� ��s������)�"]��o��C����]�*���E��n�d;��L�y��;���-4���h�X˨��@��cc �Opb=y����yb����b6�]����wo�3}��5�>�Z�j�W���i��~,�:I����	�]��UDs��$NPW�8 vim=A�ƀ�|dx<R�jY=#o���^��̲���IԐQ.�ī��O#���"��a �ˈ�i�P]/#L�]ZkK����'�:������+.�uAk(���aJ@=W-#�<$y@	�ªR臟���ch�����i}HR��2��-<2^3nf�tt����I��M��\"�}�DN�D�
����xǤmK���Q�%�|�n�����1P�&��� �a���ݪ,p�A�
��ZY��&�F�>~k�5�L��b�۴l�4:r��a��۔P��j5� e��̅9'kD��K:jjE���l�k hͣ*E��'fc�6��ICX�HLI�+&�����˭Cv6�}���*� �o�1ғ�UÅB�.z�Xm��9��ze���
���3���ϻu4�^�u���pE]��PE��y��Z}�$��=�
GF<����]4�@5��g>V86:�4�R��&Ϻ?JH�p
نӃ���?ڵ	4���e����d;��E�&w ������8`�65�;��uP�fi'�C�0z^��4s���9�2c-�J{��f����֘<�
�0�%��Qt�w,����!�J �Xk	�)&�yy�G���8P�����p�[�����%�����$�[`��ClB��m�O�7K�V̅?��G:*ZT�aЛ00�ɲu
5`�:\(1�=��W��≩ӝa�Y�·�y�`$���/��~�|������}]��!h]��v�^g( +"��+�Lq�������{6֗�:�,�-�G<~a�W)`�q�*�v�xKp�lu1�s$L��r��rr��`�����~?xO{g��&h�c�"]Q�x-K.�j�\l��'t�W��/q&���C�Uf6�6'�-ـ"��c%����a9_���ԅ�����~�v�Pb�o�� .�F[n�1�*�,-�����2��5��w��%x�l�ŚC��,unL��k?D��g����6��C�l-�9������=/�`L[Y���m[�΋����h��ګAȍ�_��%�W���d������T�����1ԟ Y�M�g�������E���S�aAn:Z�i���ղ��d���Ϯ?@�o�����Y/+gG�h�[���v�Y��HZX�#5��A����E���k6�c)����4�:сe���	9y<1�.����oy�Чs1�ъ�ބFM�qfQ�5�w�g}��P�R�6@<���ډ��a��?K�~|��<Z�*�j�zK�ͨ��E
�m��cbci0�J�t�Q@��m�ym}:��:�y#h;ٚ�4����М��+�C0+���.��3�q�����XgDc]@x��I����7�R�ߎ��Kh�%*��R�����Wվ޼`_a+{*
tbV.����V	��3���d�r+�cl��������&�3�F%:�ޙ4@�.���"q;��r��zn��@�� -�zK���Nt�z����w3� ϥ���Stc�ɱ�?�<�T���1ȗo�>k�f��͘�ׁͭ�BeP
����Yٳ%ReqH����pA��&7� Y�r^�������uMu]f3V���e��M��k�\����l�s��K %?]���zi<
M�/ 3��*#[��R�z4Di0� ������Ȩ3֎r�T���O��e谴 ���7Ԗ1�)�B"2K2�i1�w��y� ��f�YA"͖���ỉi�w�T&��XT��L3��%�6��z��`�u:�U�FJ�����e�P���x�G�"�{N@s׮���4@u����PS��p��Ĉ&%)�p����`�{�
e١��T���8w;Rj�y��bH��_QWH1�[;��s&,�x T�n�t�v�q+C3�ӑ|M����ݳ��R��P��@�6A��o�� p4���F��r��J��|�[�,a[��0n��!�B��}�|��(\q���s�:dީf�Nb�"�ϓ��`�W���[��fIΗ'D`�S������M(j���W������_Vvs��f�k�]9'}#�~@sf�IVd�@p�Kı��XCf�E�@d.:�(E�� s؇�&��]A�}���ھf�*�%"���.��}x0�W+��q4����4O|��i(P��lV�S����y���[k���g��r2H�G�|�a$+E��c,|ꃱ�,Z��B��"�E˷z���'�[�L���0S�k�B0�����z4^�4~K�i���*T�V�3r������>��7���_g�{C-���a"��������׿��V�KJ�MA��amsm~�y����v����Qw]GPVT� Q�oe�.NS.6�A��_��U�'It0w\��^	_�����ɮ�[������%[�O4����T���sy��ؗ���?i�)r�O7���>hv�LV���\���ͳ�j�����Em����*��M���y�jn[��̍]B���=;�<�)��ЬUN�`���1�������rrł���z���G��e����q�K��"V�?�s�b���%��ʅ�} �G&��9{?���z0|�^`f���p��T�.���x-]*�7o�P�؉S�ֲ���U�;:XW��9���k����!=<�������R��4|�ZXajs�O���xxh�g��1z�/||ϣ���JCU�W��D,ps��a���\�d.N}vuIi�V�JE����G2ί�V��-3t�� Ǚ]c9�a$��F����Y�꒣���E&�8 �l0	l液럽r�-�v�Ge�[�m�z��J�w���=0'����RI�n}�����ڊv��
ec��}���*@��wv��*��]K����_���1�g`}��#qFٳ��tI�3��sKU^�p��Q��J�c���M���a|�J:��C��8��6���A��i�b��U����	����b�}�\���-z�ד�QD�@B��[pT<�P��_:aB���3�����s����CF�����<@R2����r_ףδ�%QڀTV�6M�9�]a�%}��{�|�T8��Bvo�B��X��%�7�8�vD-Q;����=�z�O0�L	 �!n*n��=��]5h������O����[hp��2Cs�q������i'k��[:����屬�����n�>�z�w9����vB�>�&�_�������8���`m�)�d�� ��������}���N��m�V�'g���ٟxEF|�0Jn&�PRf�z�~բ�2}㪿������5Q�×�ͫ]�!�����8� �ٗ���.r!�Q�>i3L���M�En�B�[2�C��a�G�UP��f�=`
M���9����y��;/�����Д��B���1�i	j���kO�$�����p3��2��/��ݾ&�&��!qs�hI�ཀ'� +�������RP��IZ�+y�׀b�a��8;��j �ᬘ�L�<D�4Bn�v8��gs���y��Q����ǥ�p=g��r�d�\�>��#���w�)rO���>VV��i���J9����ҭ����Z<~L���t�~2;��7M����QљT _��:�⠻:*'�)��'a}�E����=
���[P���K������yM|�˥w`���y�<�  �8Ț9���!��D��_�$I��;�4�on��^-�OB�L��.�+4J(����,�hT��f$���wg�����w�tz�h��-�0�`���g�q_�l�x����c�v�8��u�֣3�J�L�~L��� �6���a���<Cu�.6oTU'։�e�%��$�*�EF�a�ե�11�K�=�l���Xՠ�˩	�?�kR�	>&&a��F�AN0^j;�;q{�B#�l��)ZT�o�	����΀�c� �W�*$��%N�������Đ+��xc�R�=a�i����V�ǼM�B|����z}#*l��3y��\ѯW��w���qsʄ]�����+����������������)˔m��V�b���\�QvP���4-�?�HmVp��ZA�[mvJ7�ȅ��:N�8l��D^�
}��fW2t	E�12�"E�p~պD�F{����������dZ��}q�@�"o0M�h��{o� 'M��:� ��$�@a��:��y����0  4��a�;yd��B�7�,p^���m-�i踧�XV����6�ܕ����g�jmg]��������OuO��%^����ĺ<}���tkE�P�'���ReLE��"�Mz���IN�.^h�h�����m�Q�z�B�G��>��,)�l�]��[�����M,N�V�B���������1�(���p�*��>{R}��Y��d'�r'a)���boe���_��Y��%7��/F5�&��e|�Z�_��ɔ�Ysh�U��C%[!�u�ۑ�~E�ǇI�w[�N6����a/�(�p�P�%�2��ŋBM��UFr�eI^ϗˠ�K� ��m���t(JҰ��'n.��8�]��g*vʱ��;�p����bkO������1-C���+���-jY�lY\H��ܔ�҉Z
Q��n�o"���k��ջ>{��h��� ��O��`PO��`��L 
�a~��5����<�+;��.��ipq�"4���t��p���b��0�e�̋���ζN&�O~���(C±�A�\��!BԃI�s��5�<�yOE����`#������n�ޜ&�w�ã^��Q[S.y<��=�:����fpm���+�j.dDX:�4��{�X���ϪLHD���އh#Ӷ�V�� ����e'���U&�D�W�sL�/+�ɃS�V^E�N&D�U��^�U��c��Y]��{�J.��:'a�+����a/,CCUx�ۈ��[�A���J�$�
�"���.�2A��xgz(찘�X+CI�*b�xI��#ny��T�'��᭳�T�mx�-š�(����dh0e��pw����kC�n�n��_C�򋛻9�Qcʡ��3<��HX���I*��Pn*���}p���:j���I��O�7�A�!�S�ܭ�JT����PE9���J��©p�G�j�X�����fل����T~(o��|-��DR�+GVde�@\"$<H���[_�A�bL�<�?���&,H`�MB\��� k�)��Q�E�yc�@���D��N+r��'h�{��3�8.�(��3&I�&�AID�L8��Q؈������L�쑋����陂���85c6vB1��9;��a���{*h��ӡ=��:4B\{�C����r���T���ҡ:�8`Ev�v�݃"����X�&�K_���#z���E9��|���d�OH"Y���T׉�hB���<0��2��ʞdS8%�F� >�1��HW9b�ƫ������LW"��\�)�JX��̼�Oļ0��0]��L_੾��c.���o+&pp�M��x4ţ����mD!D�EG:�T��H���և��_D��'�2<�z׷E��Y�8y����>+���x�( !v��?�Ģ⺲�C��Q����w/Nj�<ZT+^�hL�lr���%ߕX̕��������+d��z������rN���ֵxO)V#�y[cyv��|�K	N��FT��S��~4��.��GT�;=�i��E�i���2������k���o�?��S�~Q��j�e�5J��,�ý8�-�f���H���?\��PDv�&��mc��&�-JIA��;`����q�*�;NQ�e2m��=S��߮�c 㬦6����\;�TXޓb�ה�X�9J��]��o5�aI�L��n��g,�!�p%�'��2y�+���*�!�j."Gb���"#k��Ȑ�l���Nx�ᗯ����'�Lz"�D7H
#�ڡ�Z���:V;O�-A�=m�Z�|�0ч��R�Y�H�"��D��3�jIf���K�D��#�ki���z����D��H�Bĩw`�{�C��Tף?1��ą�*��ϛKur���ތ#6Ott@w�o�w^d.�����=f,o�4M�>'�'4�RjC������S���h �Q&h�R��� ;����C�V D�jOE	�i��j���K_$�d�q���v�"�P��:p�n#'��;�6r��|I�ab��b{��?K�ʑ�E�Amo�10����/u&��0r�B{�h.���xݧ���3��b��~�X���]��T��C��j�؁W��O���E����C� "��$����n��ѦC. �=�U�E��XB��Nּt��cgC�1-a.z��֕�F��� ��/���9@��V.���g:�R��>��I�.|Bӄ�.V̶�_w�g�6��ϊˊ����e�6��u���K'.*H`�q�i�#�b阛�M�-�GxI��`�|���m@�s�q�9�H-�%J|���rX+LTR��+�I)�|z��#۫r��_��U?1���/#={\��"V�'�>���nL�c-�(1��]D���gI�`�f=�7�uoI�	|!�ٰ�֮_&>��H���,^e]>+�k�b�C{�[�G��^T��ׅ��r/��'$��]}AOa��[}8͐|bv�X01D2��kF,a�:���-{���9�8 򥊵b�a��no�?� ����C�v��sj��?\&�=��@�b�߇f�#��n(W��1��J�n��_������h5Z'������H�4M(�H��_�}�D�\�-�IQ�Z#�r4�	�-C�G\�o��U��F�����%�w�Ux1�-	,Fp�=�~\�p�AGcB�u�e�"�N.<;فL���J���}۾�h��aZ����b��#�Ycҟ!i3��ڪ$�
�(�s����ǉ)	�G)-e;B�nl**�Y2�t��{oؕR/��gy�![݂���è��`��j�<�{n�M�G"������?���ۦ�N�<'�LohN�u�y3$�I	oub���E����S�=�S7���ت�޶�m�7x���2������H�3�����'�+<�5�H��(�B�C$4���9���'�Ω��!��W�U7
*5l��9e#q�k6�����z�]J��}3�TH�8�n}~Q̫�A_�8._�D����sC^�8us/c2_��#L�l �Mm�&��V�E���$�H��F�7mP_���,"�P�L��.#}�V_��&O�4`������r��CX��@��8�Ø�Ξخ�[�Yr(k�٬��(X�#�q��]A�Ĝȥ�
\�݂/�h_YWE]Ç���ٰ���2�:f���$ ��T5�t�Y�s���o<����۾���8e�_t5���P��ÿ�3ꓻ��S.9�[����2<u6#��:0��%����t�i�(�3�-b��W�W;C��8��ւ��˩�L��I<�L���[�#�"�����.�ϪÓ���9E�Tˌ�y��S��J��Ҏ�����1&�YݬȊZ��u���!�=�~T�yA��x�$z�m����R���������a�� ��b�B	net_hX	�w��1��v��'=�*ܝ��h�EP�%b��[��j���-����P�*94ql+��s�k���IX�b�T�t�ou㑠!ځu��˪؁�A�V��y���;Ԧ񡆿������,�nS��V ZӼ
��A|d�:���&xe���b9ܕ�r�[Pvp�S��6l����\�$j�Ц����0﬷�l����9n�Mu�ܣI�Υ���ݸ�i��/��&"�&�ș��;��<��S�{�O\nG�KT����qf����4s���ޑ��'���х�*�~�VN����n����41EN��v�!�E���Y�GH{���bf�4�LR,�_I�q� �#U7J�*L�Z��N�A4/����9����'�s��4s�1㚹k8x��^΁+:�x��i#"��wU���r�07��vj$�|f�R*����;<�J�d`f3;�l�zG�?����"�m�U�?JC����� (�Ym}gL9���0�n�+�\Tsa�Y��P�U���)j.3��SQP��)r�K��j�D�S��6�����s��'�쿲/A9��t���P%�"��{Ь�+o��Z;��7d?őkx������h t�tj;=���.�š��P�eS0������{2�E�γ}9�.�����(F�K@5��E^co�o�c���ζj�v*���
�`{T1�6���~�_#�dUm��۔{+�n�o3z��ph"���p��13ۡ)��C:Ɖf�x�{m��3�߄�lknu�yYtHEiq�Rz�b꧸�ч�V�y;!��ɘJ�)��o�|���,m�~Y�cF�+�G${!���Vc��oIѽE�ت�̠Z��*�(C��(�ι��$T!l}5CK7�4�pxe����.g4~�4<M�Antׄ5NL�X�\7i4+�O-jK��Ւ��p��|���Gy=C�N��#�����/H��ݿ�Fp�
�m����B=��������,���ºK�BAg!���sn�[ψ`֔'�ki}�;Y����i B�ۋ�- �)�@�n�ea�U6��Xn�xէ���W�Io�We��`����ğ��}�G�	R�TD5����D��ސ5>�ش��v5Ǝ��[��G]�D�9�B�w��y����qX��|��9?����%I�@a��$ �F��dz&���CԐj����Z�9Xs���5 J�؝m�'U1���[Ϥ���@*X�o�P�h�����x�����Qk%��E6���8^�� �!��� 8��K�V���S������t�h�Z�~����q@a+��1IԖ@m�ua���^4)iQ�U-۬<�*v7,�(F=��D�`F�D��c��+�k������1	M�@ϛ����q�e4�Z[ڰ���d�Rv
Z*�Y��@����>�zU�Y���T�U�k����Ikt>�l�[�)�����M!�Si3X��?N䩉����M�Ī�ԃp������E��T!e�<f8/�[�x[l4ʋ�[=E�ފK6P&�������Uen�5&&������|�D����Q�-�A�ӵL�n�� �1 ��ȚRH��e��f�p�h��mx�=�m.���Ts3�:|�	hm��+��
j����S��*��j�{�ZS�
q}�Y�1��%�ȯ�29 i�M
���9&Z�6|��<�j���	�O�t��o={[04�Ra��
��Vu�('���X�����+��
2����:���J�V7��Ut��Ю9���(\~�jA��tf7�NtA[�i�t��$���B=���ႉ���*� H(�k���	�?��=�v8�EO��E����S��dS��չt��'(H�nuq�6���G�9��P=�8�):�����I}���#�.fF�&�F�@��~R��<��������~L���#�Z2�4���C�F�T�;6G^���A/�a�>��	ʀ��0X�zI,�CҪ�IB�.���L᳟��v3E�:!�ˆ�_a���K�Of���#���le�93�)��{T��~���V�/=mj��0?�}��Wcg�;-]I7�+�J��F��놨���`V㕿��=�5�m�y:���^���y��>ף:3��Bp�?�����������L���@��-���Z}n��UϜ�"-�,��Qn�S���uy�~�6���������^0����x��3j�s��~�5K!����l�����9�	�2FK2�~V5����@BS�2b���Dz�#�������Iu�mY?9����v�/Z�>��io w���]"���r�胍�h{�[�yIe���'�`<��l���۳���&���l�BBۄ1z׈�\;A�J��c�M�;vR��B�2��hr/��h����9'Z�ķb����IL�W��ˮ�&�`�IN4�IVȼDb�v����Rߢ�Z�p�f[qݯ�0lNӤ��!�1�~ߒ�h�7^D�Q�?\�_*�����0�$F��*.��r���J�2ה\�%��Xۻf˷�������)�Ԗ"rU�������[�f���L�E;�Cئ<�,�
~�&�{�*��Hw��5|�Lr9��U3'��ґ>�C���/a��y^]�gǨ�90j4�eP4E����s��m������av�fAE���X %���@)���]�Xy/����֕�Uw��C�r�LT�VJ�i)w�Zd�ycձu*�tC�N���eh���Ky.�oFo�g�E_�w���c�<��cp|s���"`*b�{��&�CP�S��Y�/� �Mw�'	;�<�NAO�BE@
�vM͒]~��^����ڔ��r���;�-�����&��Z��"�E��r�#Z��\G���a��bE�?k�ޗb]��Px����s�^��ڪ�}:���{��q���Ƴ9µ����ˢNn22�*Cf.K��Qa?�9�-*��>���N:�Ɩ��X<�����`�+-��.�kd���Nm��B���j��5b�zL]�K�`�c;�n?�]ޡ�EByG�=3���XpPλ�=��Gc�&e�<N�X����!�BP�ܾx��k��ܘ�ߘ�ȿ���o�ɷS)�P��������W+�l^��O����^w�܋�� ���su��GXGIe�������v�Й�Ⱦ�e6��S�2����w�<����;�xyyt?y�� k�,��ø�����(�/e��!��v.��E�7#��Z��|�7��
�;J�I�ä�[I�OI�{�к��>}��2~K]��{��<�1@��bV���$��r�S��K�y�j���N����u��1Jc��|F��p�ޝ����0�#�р<"�e�jZ�d��I�{�疟;�FVhsg���+�پ�JI�U3�J�H,dæ7Dd'��2ӫ=�"8XV��6�M��5�CҊ���
~���Fy��`�����|8L��ѓI'�g"U��7f�İ���*"��P���C��^�e�mw�6�@��3"�f7r��h&D\�#ƩqS��HB���l2|�|<XQ'������S~�+�n������Sq�<w�%y����
B;崙i	��`nm|�m��g�LpK&�X3�*[�9��u��MA�5�)��we��
��-��8�����Rభ7�{�{ª�;q��;�,�"Qe�����Mz��`�af����{7A9�� 7�0�P��ڂ����#��7���]0�,R9"�g8�`�î�=�����i�)���'�v�V�Hv��N�b(��Y����L�x*���%���d��f���� dBӍ�\q|�М1m!10F��h��U*���i|?��ϙU��U�档�K�p���%���)���N��,�a�Շ�<��`�o��jt�p�@T�Hv��CQ��Ρ�@D�AS%�/Ӷ���̴�����l�0����׍��+��;c�|A�>��o���cS|��a6����8���P�"h�	c�tI�q�ۙ��N׳b��Z�t.sq��7{���mXSZ���I}/m,�(4Z�1{�gpf\6P$��f���@VNb����<��*'�����Q)|ׄ�Ӭ�y+A��Zd�4)�gU=�r�=;
��^�7���,=ҏF���}�ɲ\�\�iR��R�P\�@_,�qඑ�CǼ��ɲ�En�1C:��>s�Uϰ�g]��.5���E��Z�r�"�,m]6����@%�c�I��@Pͫ-��Y:�;�m�hD&��{_�ik��[����q���F��<�JR�ړih�vCk�����cv��h� :��n�����T�Wn�E��_��o|��O"?�*hp��:-�T���N�]:��u��6L�ۀl�#��4�s�ޖ@��?�vR�5��{)KI�?6��_����:��H�\���[�8!~�֪�Qٍ��0�*ڟL����V
ͭ��]�d���5}��T���>$=>.��bS|�����3弥��.�QY-��^nƒ���! ! D,��9�}'�65�Z ~�yՕ�Ԣ9��^R=%f��m�h�h]���He��U��䜏 ��$J��_�*�����'�����g���)BU̍���Tc3�w�H�L&[�*DS�w��Q�"2�� "��̫ru���#׌fW��w(I��\%��OY�Y���/�w\��P���!o	^�|�fq��iSb�NVKv�G��#�Æ�x�~�˘x�u��%�����F�:&�k�Z@_�2NٿA�]t/�Q2(B�2��~~R�i��?�P���bFHI���-�� �C����<M��N�}�p�xaI���f%̖;�gT�]�ez���m|7���r�|8�E<��gi��EL#Ωpc�bt�]:�FՓ<Ҳﵦ����Ԋ݅IM .w	��
La�󐶂B��L�� ����LP�]eǹ�A�����X��/�r�9G��n,f�-�'�������R����v���AG��4q��.�P@s�F⺡��|
+����0}<�8;r�D&��Y]D�G�:x���<���4�;{7Pv[	\V��j��b�KG����)k�$���Ϋ莃;�##����S�=d���]K&+k��K�["Vw�;�I�y�fW��B��m!�8I�E�D���w�n��w���7�A�z��fƢiHO���$L��Hs��nr��Z	}]��Kb��N���S?�O墅�;Z������;��|�i�N]�������H�=�HT�l��l�E�}�d��1P�1��E��k���K`�x�Ǡr��iJ�1N]����xO���!j-���|%��e��E������a`����U9g��9#͝��牌���U��D���C�Is}�-���)7��#^P"�8ˌ��*��k@��>� ��#�7��s(@���4����M�Ŗ��خ�}-F��sO9�R"=�C6�;�TUY�������ǉ}���	���&�̀�Ҭ/�s�4���q��<�H���V�Y͆��ML.�	��H
4�Y�>���b���I�1��b�kȃ�������y\��YD8��Z��!�aUM�����s�j����Hn�Q��j�
�|�Ll��J���#^�7��[�M�3E�Z��k�y����js`�< �wn��J�ao��oX�}4�הB�=u<��1c��&=�F�@�F!c�����2R\K�<\s����J֩�\����RO��+C�ƜC�Y>�{2�&Y��{{���_�f��m5�i�Z>h�)gC^b�o�]��3#̘l��
��nW�o����@�oc("�%��wg�&���F�7�d�,�
-Z�=a��B%��rJ��As�$��Ը��!���rA�')��bJaŌ���4����+�ij�qMF߬Dr^S��X���Sx��/��%��G�{�<!~u��P��Ł�V̘~I��!4SI�5y�h>�J�*��f(����S��u�/�`�<���Dv��̃.J���_�?C،%d��X��/��jG�f��K�-g�F׊v��\EgCj�t��PM~��wO�i�<^a��E�r�7�Flpǐ�A���U��N�#Ax`�
H�5��Ӝ����?+��I���ؗ���T1������v}�0u>n�P�\��\e1��O�9ny��ЬW~�X:am�)��ɘ�f-4{yΰ���"�t��&#<�:�`(�}|?�0QeC$f]��$*���8Vt�Jk,�����;I��ό��#�����]�`�6��=%oh���qk���5��X;9�$�"D�7�W���W'd��r�H�sv=�$'�ޡ��e��JσF3�8<�ɎԨ�1R�_y��_������U<�/�Ɋ`��x1$9׮�_�:�#Z3�NyነX4���S�ZOC��L.���t,:;_��Myer�6F�d{}.��?x!����M*��e'�b=�f��a)����2��}=�U�H���v�B���XO3���O��7$Z
(&����ÙI1��^��W&�P�S�s���zVn�����5SQE�3Keg.Pk�$�������G��O?��E����m��S�N��C�`U���Qq��ܨr�{��PAd���%}H<�S�_y,W�q�X�tJ���v/;r�m��D������V��S�]a�wb63�E�|�����W73�f�̘>*방	�Sؽ��vd�J"��Y��@�c�!��*�%g���^M�_cV�.=�?�v�;y�^�By������)�Q[��o�ph.	&�����Z\���x�����G��]u �$�y$�Ă�Re�I�.Q-����0��i�d��RUY`���O�"ٍ��<є�;�5]�PP�,B���_�=C.��f�'���������gۇ�$��(�}��񤏰�Y6%�W$-�^���ߍ���HS�}�Q��D�g��L�r7� ��_n���� �z��L��;��t�vϹA��:U�����I2��J��5Nɦ�@_��%��k�Iq�쥦Ip�߇d �5|��N����Vqp�/���a׎FaƎ��7��}S�O(Y���p�)�'�p����L[�9Â^��}���w#1��@�����Q��ԧ���~�M��;�����44Cl�6,�H�??�b���q��)j����K��m��T��E�ې��r���ި�)RP����_8�=����v��U�"D|=xVU��X*�h���B`��ק�"�&_ XR�'����
��v�ٛ�����WqY����q�a���fȔ�����_[����� U#�!��5r��I��5@�������,=j:3�A�Fo��g�DR�==/ϽK����m������C}
�m�U�d̶�_Q���5��l`n������,.����g.������y�v�]�)�a���	R��~e1_�,��o�1)]�@�G,`���R��<��`����ї՚��1��ڎ
�h/S
&��_�2���`6�D�8{�;X�"ٛn�LT�f���e+T��'%{����cN��m�\�2���d�F��6���P��{�7���w�`a������z���͘�2�j@�X�������oF�7�)��q�i�:w����W�'�Ì[t0~s'�_��>�e���G��^���hg�K��~ ��o۽űF��Y~�v�.`q|c��?�"|88��W�f(��"��5���I��-S�� �~�W�)��GI��z������3��G��!��tL�Z9[��J�;���Ї�F,l�-���/���M����.!>��j��!�(��@���i�LA!;#�l��rH�1Z�����*d�Z�ƃ]���0e )�s.��2*a7�߷�R���27uv�b]QټFdR�RdB�q�Y5���HQ�灎&#�~�0��E� 2���&VY����?Ƴ�M*_��\�!���TfޭOwn�K�R��;.�+ͅ�Z�%z���)�ta�Ѭ���M��^��}�D�j0�Ƅ�H�{��g�zb���̧Lf���k{�͉��9�@{������?�R{Ӡ�p�i�1���-zn �w#�_E�Ⱦ.;��Ҟ6�s����@�t���}y�� �d�&tL��Vg"��`�7�;��ݝd-�R�tx:GF �=J��!'	�w�!�N-�o����Pn��v5 ��l-��\$�ZkrW"4�����.����?WԴ4���R��ЪW��;�	ce��z����Z�X�x �6��u��_��s�iѽD<�5��j���)9�C__R�?�H^��Ѳ��Iz��7��h�e#�o����ԯ���u=�$�G
�����p���쓩�Ih�ݤ�������k�z�}�����8�buI��Z��[�e�JuWx+�����߯��z6s�"p�R3)�z�c4�%M�n�u�F��Tl��;QB�f4�D��=[W�P�X���N"����JJ�MO�ʅ�աt!�Y���Qe"��ۯ��0����m'P�=���d�\�sg���/�(�]���X㨓�e*�0體X@\�v]Z�J9XbZ_������G���."��W�<q�-hD4����[�k4}oD�#�B`� �_����$	I���o�N ���\�Gn��-G�3�s�����)�8]*,BjE�0o�O��U%��˯�ZnLENSi%I��z$�C"���%���$;ʩ����ό63~/�V���8�#��M�ζ��j�uAx9��xK�8�1�9�!�'�}�&ZGc�e���,.p:]���Q��a�#��`�%&T��:$t# �hW�#��+�9��0�/�=�/?
M��y���J�%�D�4�~�#o�o8̰��M_�V����I>¯�c�?��+���黈���F�EԶ+An�n��B�ą��l'8#��k��	`Q!0�+ty��t���eVHv��o����"A���8��[�v���`Z��J8<�kJ�b�����P�S���"=p�8�^��C�ۂ��Zb:r�+sNn���J؜̶HI��]�Yy��/�0�:��nE���.�)�rT�L[P�����f�����4�]Aۧ�<��w��۱���yV�\����X|���9����e�:�
V���8��կ�M�R�I� �} \lP�v�,wH�܂�8��ο�_ϰ	�9�_'�$X<�ʒn������M�[&>y{zf��O�7���:��$�M޽$�x.O<)���L&����_�~�&r��� �(hOSU]:��!E1vՀ�Ն��׷n�����ê��_���{�8j�yȘ�46�9)=7'CR���Y�p��w( ҩ���^��ԭ�ܰ�7.�x�"Y�c�VA�����X���j��(�jP����<�i6��Q]9_���t�!:o�i�SP1��~��1r=�Ti���A������g<��g;���]
��w_`3(~V�IZ:��IB=�n$���<n�G�۝A����h@�;pI��}�|�}4NyDD�;ƹ.)��#� m=Նw�Gʟ�<)8�­�:H��8�Y\�����u�>1M��F3��-�)td�qSNk�^M�$��醝�Q5��w�,��.@M���ۓeEH���tN�;{�C�R�#Ko*����@��E�#(�`�WMΎ9^��9і������|��[�^4S*`{z��eo� ������$�%���5�l��`�o�nA��D��hx�p]�fP��,�ii\f4uil 9gƨ�h��d�2+�{���*��}}��[��.���"3�.�{Q1��K�CWGO�'���85o���%����+p�[Dl���������$.�KJ�+]��C��3?���l�8O����.�3��L�f���r�2�钜"YӨ�:}�CD��E��-Sȁ#��c�Ǭ�����J��zEZ��#���I�:�ܣ��@�&���Zdl��T��D^���N~�E���%-)��c_x��p��S(n~�{����P.��Hjy�ȷN�$t1*��P}�G y����0��x|�Ŗ�M�yϽ����O�2G�Hi�n���h`J�}%_�b>c���ߙ.J�C����݇I�������ķ*[*�Hu=Q��a)�q)�g�kJa�H�Ŕ�e謒ŒXU��H��\Y�`�!θ�j���WզuO�6(����;I�_h���n�hG�L]�X4gR��น�����E�"#��g�mU�k&4�c�s�p6���UXӐ��V���+ܡ�GS>�dv!�x.9�k���2M�X�"��bi6[�06��t-Q�B�؂��υ�$���q�%H(vǾy&à u�V.uYE�uF����*ݗ Ԝ�:x@���n4k��~��w�*�rA��\��U�i����[�f:��H81�N:�F�I� I,�	m�i��&�x�K� ���t��0*��V�J6̠JQA�Ad;[?��=qT� _�[W7�@�Йaek_lQs��
P�uE�ќe���FP�f�� ��n�0��Q�_��3��c���Z�
o\�t>O�
{VEoŪ��.�|!Lۖ���`YJe���VsyؿA{w����a�/�;a�jǀ�<lN�LN�7�cc�ΌqU*�Eo��U����B��w�s��̰/��?N�ݐ����|�p(1l�O�J�q�Bρ�3�0r/AV�<S�x�h�������MH� �;*���^*mE8 �+��1��coD8�z�zWn�ܻ�7���O��T6=�~X�`�yz�q���%���y�sC4����)��$�e�j�6�i��A#�����W���5��Xw; .��O��:�=�7}�>� >�����^��4�T���U`:�§,��\��s�J�8j��-�i[v5I."QQ�M\^��R�|�}y̿�i���9F���yEs��� 6wu㙁a��WO��X���G"�¬\R޷�*^�'(�ۤ;<��Ж�P��󕽼��V/�N������T�tF�0�aR}3��iz�~�`r��O��'?r^�P:��"�vHV�����T���m��,�I�Ѯ�1�Sʇ(�������j��s����j���syb���R17�U��-؊Pk��cH�ܭ�a�� �'��jP�&I���'�����!�=�4�H+\R6���傿�[�Q����L�� �Ok��ߝMv�n�㾿oƪK󜌚�7�_M\�41���Y��HLx�H��ʹ���$���K�[s������>�B9㾭6
��N���~ ���W%'l)4����)���H��\I��t����s�Q��C֑�A�/!��>�W�
ꨣ����.���D����@U|��,׃1\*�����_=709ش'�u�i��g��Ƶ^.dL�^���?*�Z��[����F�hM�eِG��z�\4���@G��B����y0���n$�҂sa�[a�H�T�`�_���
��&g�fnn���T���;�Ό�8����v	�@�J� `vTБ?bR�|�4k�e}sY)� K�����|�"45�5:��nDA�7Z	|�$���	?�>��-P|����c��2dY�x"SyX
� ��Ǳ��s��.���v�[�j���"�Z��8�/�XY�t��y�a!����Z��l��ÊL��䊍��������`,k?��������ϓFӽ#a�>Lشt�B9������T-�;'�S���赂~Z�@�+�F\�w?^��X�Dc�u(0ul�S*kT�R������]?���Kb�^�`͈褛���kBR���sB�|�豀�i+
d3��UUwx�+�����s���^p�}H
ŊL��Ͷ����!�%�9�l�C�1�g�������C���+���m�t7?��-}Ѹ�+�R�Χ�-�R?���l�q��a���ݡ ���j��Ӓ��~{��*��;���ERH����rDFT�n��`o#�6ܛVz����`��}c�"J	���a�O�t�����뿫�U�Jk�ޮ֦�g��}��JJ����y+#���M �{˂�s�_�D�c"@@���xG��R�d�!p������q@^ZJQ&�6M�J+K��D���AZ"�p�5K��K�Y2�N��(k���C����z{|5'����T5�<\@l8�j�hrS�V�p|��i�2����R ������[u>���r��k?��X���������o#t��Pv:b{�����I#�K߭Nx{ô8@u��&*O�%t�S�����\�����][ӨjS��"� �Jvl�$�m)7@�����z+��y��U~E��p�P��{��ł��*�q*���6'��t��2��"m]_���b�b�f��h�U��y��*��:S���?�n�	d	�FqM�j>���u	���lV4 	��N�b>c%����"CM:bqDo��i��$�~k;*�rt:A�sv����,�x�@�V��.�[X���L��ˤs�s~�ud������_�C��>ըEi��� �Q�.�IVˤ,��o.�����8����x�l|���F�d�uDb��w�46�U��Ju������O��-� p�ܫ�0����	���%���gX�%R�a��W]��^���]�p	��+ɒ����u��'!k.Bօ�2)����h�OZ�Tmϟ�(�L�t�����k5h������BԞ��F8P<p�1�$���[z]X�Q��i��.���B$gv��m��@�r쿃@$�ߤ��+67������^��x���ûª2Z>�F��6M�
˰��0Eog�[9|Z��O����$7�cI��\2ʏ�=*`*q7ڻ@>Z�hW���5�Q�-����\m��Yl��Q�I��}0�~T$Ic��U�H�pxi/[;�,��8"�������A�]��)K���6,��2@��V��`��^RdNud]S�4ծt���4��嚢|���},�U��30�E�_��$��3!�CjX野˜�]��-Ԉ��{H�T$ 9�D�^�-e�yGᙰS+�O��zm���RκT��R��B�:�ł��*
�LL1��l8��o��_d����+�8^�v���.���+b�w�I�Uv}���_|Hr���.�xw���̷��r��w�w�Ƽ�?{V�� >��1}�ʀv�;�C��~���3X"���1�����6�@��+������@SA������G�%��J�K�v�nE����� ��`�z��.Z�J=7?ĝ'I���G�oE?zi�%����ԇ�����@��辉��T��Q�((�#;z�+v$���о�}4���Q����x�Y�8a`<ǣgi��\���W(���d��g����5r(�u�^��1!�C�#P�b�qx|��pO�uψ{ͪD�?5	�"1� R�ݏؒy�G7�'Cek�j�R�bbd��qa���o嫭����~���r���nvR�<n��L�X��Q��(N�_*(Ϩ���Z�Lr�fLr۩�@����4;��&��Qj0�h>������F��k(7]��{�RD|�I
=%��(��G�d�ݟ
�h�>vA���x�5�2j�*D���@J �7m��(�H�:a�3o�<�B'奈��	�D��	4�KS\��*�Z7\.��NSq��)6��("??Ӡ ~��L_�\�mH4����1wl��� ��C�Y{.���\)��4vh�栏�^ ��C��q��?^;�[��\�J�n�<.3H4{��;)�q$.�ۚb����s�L͘e$�8��dKf�ԆU"�`�^�&������9��j#�}F��^$���R*?qe�S����p^Y�Dsw������*�𤌮� ��*6��q��I%�Dy| ĸn��j��W�e3�ѥ���O�bKOx;�{��I�(�wB�h�~J�¡�.�끳j�q��\�<�,�=uzJ�5�u��@)Q@�P�5hK��_�����x��ja�7P��'�������pyr<m/~7-����xb-%���L�볞yl�U��|�OV9���@gi?���i�<�7��V4�hM{����M��-n\����tW���*>N�烕a���w�[����Z&-(��"O`���H��rȸ,��������|�9�i�lލ�+�m6U��j쵔G)�FYZ����7�T	����*KhM^��R9��ɝsInS���>��.��伩Q��	@(��q��Fi�&<Y�uKW.Nv8�v���$T�dB |��Er��q���&�Z%ϱ���|�l.�|=�#UB��"�f�R|�A'�C�k�O��;��$�S�d0�Vr�-�΢�(�� ��I2�.=_�o�^z�h�Zn�>�{�p���t_m
���|S�b�U]�J����^�t�v��"(����z&�0ɚ�C��SӅ򬶧k�Tɛ<�u��ᤆ�G%4 	οБY�̖й�k���<Ҏ��[��z��&�F)�nå�݌͉������3�����A�gp�zJ��e13��wJ�S,	�RKn��ܖ�_<q��	�]k�;J�L��H�3;�	R"�ЦzS+��?����u���Ӓ�yU|kDL�݁b���FX���S$eL �\6q���G��4�=��?SD��W���X�ЄQP�Z���Q�C��U~^���Ԝ�z]��E/���P|�Wè|<P��$)�)�j|љqn@*�Z�)<}:��+�/[;�H�~\ŗn���m�������Ck�8Є�E��o�џī�c�zv�{�c$/�Et�QmR�--@4�aKo\��߂�uLL�u�-qq�[!�7�Ǻ��FC ��L�!
,	>�K�`
��pO�4��>�V��3�-��]±��uϚb����?����A��Ь�j�:�p��8G�xSYQ�b���k��z��05(���S;)����� �����Q3%'%:K���_D�&�]�1��	0�Y?���k�������u���d��c�0 {�}�x�X�k^.�7V���q1�؁�%p����!-�b��j^�����kb���9�P/}��I]�W���'�Q���o�Ⱦ}�{~�0������9/�[zr�oN�������0�hmD}�"�j��^���� �sk�v#��n��i}ѕ�D�K�}�6ia|V�ϛ��"�Q�u2�p��	B��O L���
^u����9��&el�	¿Ep���nJ�/@�M]�
2FR��V�����\&�߱�0;p�{��<�M��H�`�X��,/�Y�r�)I!oP$i}�C O:���q�L�q��r��h��D�j����{�?��Q���e�~�]Xs�w<Q�섢-(KЄ���#d�f�R�=�BxBj+GI3�a;vs�Ic�Do�ep\�x��x��Axϋ U��*(Ug��-v^hZc��Ϥ�З���s�58
Ҝ�pX�'ŰP�C)^��W+;(�Rp���?�Lf���Z=O�����6��)��5���U����Q�����t��[W��6�\�����:p�6��6Ub�K��c+�Rh���$��T�Q�'%ֻ�)��|&©�pH�藥�PΨ�B255F��bD�Z��$-/�HO22lI6/;RN�� ��(*%�N_�H����bA���� �� uL֠�n�'p���gQ�����
�5n�a��
�����'�h�5# t^T�p��W?0�D��;�;�S+��ا,�L�ݒ'�ʥb<�����k��4j~
��}��D�������o
HlT��\
C�|�
?�5:�����k�}B�`�a����F�?�/�����������v�^v� ��,&�B��y���b�2y)�n7� �W��Yl.����5^�<H�|tD�C��[�]f
(�0���.�|:���[a�4:��-��0]jZ�wڠx�� ���H��*��y�<J&v8u����e����3_��)�����N�	��uxz֫�Ms�s����VG�33s7PFv=�A �t~m��lrDH=���^��~�l�k9�ULy�W��鬇"�uq �/��1�2��N�����,�J΄G��z$ڽ U��BNTs�� �Q�,]����1��.���2I"�$�X��Re�X�~�.Us�E�UÐ�[|��.fNo,�tʔK��H�M�_�R>(a��Ǽ�������k��KZ}$����w��ڎ{bJ�Z�N�� �p\��h)la�/��Q�����~F6I������\�������ɀ�T�R׃�g*隔d(�U�`D������6_J��Z��CضH��\���'-�����3HAM�D�	��� ����}b!�U�z���yr(��?�A�O���X~W�d;���J�M~��*
�dU�t��¶��,��0���@��"$���>��gC�xo�uo~��(x\����cC��J<����k fJ$>��v� #�z��:g��|�M�.�M!�Jl��-X96Џ���([��bZd1"���қ�ʼ�qUd��1��}����.T,a�L�K6��?�έQ疤���mr�D59�c=ԙ2aNÐ�.��\�>�ߛs��p��;
�'�+;�%�2R��x��J�D�g\���o;2/����1�p��.��4�i�;���Ԅʫ؈�K!x�Ĕ���̭����]v#C��E^���>�{"5�;򮹄��ߖ�熁��S�E�ۑ� r |�b����WƤC�6�a-��	��B��/������ɩߚC
��u�T�d�}��a����W� q�"ry����}���Rp0��E���Qer�{IU���TB����ia�Ы7
�E��UKS��g��yw�+��X(��(��d^�t��8�}���?�*-�^����Db����ng�E6/�$�7R�2Xځb����D"U�8�,�5u&ְn-A6}�j��2�Lx�qȣ!ml�kR�6+��5��]D���h�q*�a��O����hf����RL������Fp���F�r�gQ�6���k`�ևzׯEN�C˕�i�EF���u6-kc1���<���,|��G���,~�\��(�Ov�x� d�֪���WFwJ�����f��PjK=<�ȟ��Q&�J���? "��UN��/v����Q�����s�ˌ�V��ov��Ƨ{7]O11��ݹ;�2�LG�|�����ZNǤ��y�`�&}�������)m�̲v�C}��CGɏ��$8Ʈ)h�LДQ��)7$_��(M#AY�#IIb���Wx���ۀ2bM�[�ߜ/��G;V6��S�t��1�Ͼ_HRi���3>C�%ߍ0m>nK�-��K辖f�_��������P�ՔX�F-�|/1��� ,�ٜ,\�㈏�!�R�xѣlV��<M�~��t�M7O2�X]��;F}f�в������i��?�4F��]�'�R����b��$qA�F�.���3�x-z�B1V�˚χ���\��4�}�U�ڤ��#��^����p ��t���*`Eq�w~d�����`?E����j�'-�%�Iy���*�7	��`�A��퓽�36��Of�2N{z��&�՝��5�tY�.k\����VIۆӛ����$+'ZD��\V�Pj�O�ಔ�̪?�
Z�p����VR(�T�`k���+؂Ya7��jv�<��R�񽚾vGP��������!B����dl��|�>Sn�s�6pB��F����~{�)�𳃭X��2��+��$ժL��mח)�2��(W�;�_g&:9�`|�Ӌ�U���ͤ��6[xl��, O��f�A0#KBi�+<)!�ߥ�@��:@�м�S��?��҄����\P�K�+�;}?[���Y��5q}�j�Zl�:�;'4�|�+J?�]-�j��0��������Ί|I����]�mfS�����	acׄ4H1<��A!��o�}J�&��j�%��������(����H�������&Z����5����� ��/c���p�1���*4(D%#e��C���z�g|��\JT*����F�Q�����D��ė,��4t&�^�0�v��Zu ���k��d�ͥ�x�(@�m�\�'�)Cȃ��o%Ҋ�v8Q���ZP1*�M�BF{�%�~����v�z�M�SrK�o����;<�t�ު��:,~+��0Aw�%�zP�=c6���e.QC$/8�u��]i��=2e�6p�r|IB�0����|�ۑ���(��ke�����*yVH2�X}�젅F+�ظ�X	�D�����H\�m�o�c�)���!��W�f�U��F�d���`�o�E�jD���`�-���2�
zD����ZWj���]��>��StN����͈��"�k���?�/aȸ
]4m(���ګZ�e�$N@�d7sȰJ$?���b�6�p��X�2�ɪHHbE�����*�~��iC��;#V����R�XW����1��w+�K�j���f3�|vZV��.�mG�1!�#�������9� G|9k�ˁ��
Ə�E�Wv�었<��� ����EN�ٷ\� +�9F��i��Z:m������`_�ܓM�>SFЪ׷���8���������M�L"�}n'b>�W�AD�%}�Ѥ,�����'�� ��Ye�(ݐ�)�=�x0"l��>V@���񂹩 Q�Un|��gK��A�#��M$��e� �F1�x9j���f�ڜ-)��A��z8�5ƕ�u�9�����M���+�����F��4qYU,���pq���S�,��5T�oR���r��˓f�ӳ�O>&&�k�S5E_B@c@:\<^$`[�����*��ȼ�_,� �7�p)o���@(,g����kX��|��|���2mbS��A�)�qQ�%�WE��E��ωD�#L���1!�ʉ�a���n7^�b�sj�ʇ�?Ƒ��c�.� �t^~��{#�w�#�$��=���vt�s� F����A������l���ȏ���5��^��*�f!v��oBi��H��?�����^?z�e2�zN�dܟ{R��̏vl!���G�J)P�v�w�]6OמW�(����r�~��享�;Ϩ�?��Ѕ^�lU]��fl��e�Is�X�D1�e�v-j��a>�[�tw�ϜR��Gul��P��2gɓ�`Vu76=�Q�rB0�C��Ҧ���n�`G�n�&�#Z&�LC�&9�Qˀ��t��)<,!�{�#�H�`9��Az����m|��� *S�����3�d@S�lΪ���E��$o�(��K ��	�e.+�����^��\[�7�@��WY��ՏKXm8��h�(��=[���l��ʿ�ƒ7��A�Xb��߈��	�T�r��C$QS�!&�gj��N�Љ]��a�~��O�Z�Rܙˤ�A>�-��������j	HB��4Z�Y�y�h
�©�j(�15�#aL%ْ���0�`�x��%j5J�&�Y2�5��)��0
q�$l6��дDY�>03�dh���������8ȃy����!�R�ww2�?�4�W�ZX����A<�������+��p��>�[F�5�����P�	��T}��	l�-��v��|}*(�߂�����/&KW�A�O:+����꯽33B�k�B?w`��}�w���"5 Ю����F����{�w,U���q6��1��sj�� P�[T���J�]���W
G�
���c�:xrf۵j�ف%� `8�/�p�N"n��޽��f�Q=���CA\'�
k��麏���{�(�7�J�A�dS�V�+ooe�t��Bg�SN�SZ�A@�:�R^ԉ��EnÆOG�t��`��y	��RR�lIl���nJ�R�	s�Z���=��F?V?���lx�̠u�6�t�W������_YK1u���C�\|�d
�|�c��g9j~<J�7L�v ��k��fm�Z��sJ���+����fp!/G��2�c�g��-$�%��y�5��j3E�;�5 ������4��Ɯ��r�&�P�9���<��tm)d�?@���,W�&'���� u	��&Je�}&yDү�A$&=�F`?�a~�n^V��Zd[���Is�5�d�'��JK�3�t<�"�1��2����rX� ��T:C���Ǆ�þU�Sh�&=#�����V�w)���z+�o\D�x��H�f�Y���9~��Z�G��4D��~s�	q$,w�Ub�:�0"���m~U��i0p�I�����>�nWn�_��d��hPE�N<�^�쨤"��<˶ҧ�*�""I݌�zr��]�V����^?1�F������}�P�s�y����h?�����T�ZWOѤ�O�d�����A��Ft/�)�[8����%��DVYhϩ��
]�)��/+�zX�2.���zQ�ߧ_O�ّ�)��!˟���xQwQ2� �0}Tw?bH�eN��4������S��Ӥ�Į�P3��굮�Y�h��ʋ���1?K&bT?���X�f~��W�`H�X1����'�<��yMR��P`�3x���3�L8��x:������\^95ħ%�Q����:���'C���>p�4nɹT��smr���S���w���x8��e��X"�M<�0�F-񁦃�-���]<륗C�OK�b�йpÛ�g�q`������3�Z1<�w>j:.�H����~�GQ�>~DįYk�ڎ>�y� h~gR	�����(~�pma\a�P�]����n_i_��:�M����844�3�fe��F������b����hm�׆�.م�42}��A� �Y�u�XJ��s��ڬo�8�gm��փV����in� �g��6���/<F%ܭǩ��0j����B�ZmZ�zA	^���9�u��馓�|7�A�ZǨ�Ɨ6�KZ-,�Yf�^Z�9 ��ܹ"��K��B�"S�tء�T��=�2}K�aL��I������,�6h֢�{B��:%q5E;f;���˔���9D�?
;"f�2�憛����V�.S%0U��d��k���� �4>�OrZ]��gʔg�E�\�7�>f���c��Cgd���z�^K���I�;�Z�y�K}Ĭʣ����Mk�xh,�hǽ�O-!(�zj����W��F�pC���f��G�j׵��Fk���Zb���+�7��3	1���-	^5�x�K߭�&I�.BJ�.-��.i�C	�D5�G��N}��R�\���G��@F�[�֫��k6�������@$������a	��"���ZW� �u>���*�ۈ���-U%��2C�&!-0H�-��{G]A��r |$�ԉ�v��\�������y='�&�!v݁!%���T�ٴ=�"Ϋ�:_G���iMp�#/iS��P�����uP��uD�t�<��k�5�Y�R�"+�ֹs��T�]q����$�����lA�V��?X��2)�e'��]_��+=�� K�n�o��k�e��9������OuwQ�jԉX���uW�!�[�[��=��g������s�~���l���$-(i�B�(
n��K��ON%���}R�4�I��l���wE���=D��-JL�B�"�Y��Jx�p8�ߎgʈe�������i&2���	�j�\@9J���`����`ZeҬ�Ew�Lzi*��L5��~R	$G�N�{��� ��u�x� np�$��c�~��
���� Xז���&��6�?ѷw�0`�-Z�`y�'xmpRg�49M#w{l�%�y��i�m���!#�E)FEr���ݠ~E������Th|O2��<�Pmci��OR#5?IA3�(jqQ�(~��7~�������������d,�Q#�6��#���nS���`�Al/��#Ar�$�_�p���'�_�_ǅ]|r��Kt�hݟ(�x�	k�i`��ѷa0�=2�F�y,ǲn�w+t?��Vܗ�;��z��[y���q`����8�[�Bld�ƌ�*��_�J'>����(�� ����v��6�![��#A��ڞP�X�R@��L��)@��q���օ��8� ��`�Q��������={.�Z�Ή���27��iȉ��٫9N��$P�gD��`;��0X02�����tW�I��iS�!,�j���G)���*�6Hqtw7ԍ���Gg�r�0�=�!�A��u�jk�q�7�遗�X�(ԉ1`utR��	H+�ʻkmô�0Ԋ텓ܽg�z����	S+�R�nL���l^@��=�L��D�-�Rg]ƻ�����?Q{�x�.:zt�+G�TM�4��tF,Z��l���=Im�{�=��fp,VDgH�/�U�j�?zg=Mzc��桥��r���li�tv�X� ��m�t���w�����䬟��R�J�e����mF;�u�p�;�Q2SI�k���n����'_�
��:���c�7HG7�g�q����%ϟwC�'�ڱ%ge?��t��wՙ�|N�A�j�9��_�3[]e��cր
�E����4��H�&؍	����B����W���̱|5���ƞ�!$k��Tp֨��@�۷c�S�&f@���1Wr�t�]b�L�P�����^��|Gk����� ��+>"j<�t*�s��r��&L�G��fC�"�7��!�Jb;�����V�Ia�d�3�T^�dn�o�����'ǔ2aйErTaH��n4����M�3"��4�-�ɻ�/���1��k*���IK�� e���(m�S7%�����ہ�������ǔ��*�������»�����g_Ig�=��u�x�t�OyM��Z/����^��nZ�rMn�#�x��|���\'[/���PL8�UbX��!h���Ww����)�C'46E��Js�ft�W�	�*?�b?%m-}��s�$#C�B�H>ȑ�����H���騪A���H��#A�~{?�*��/)F�I�PG������̐��B�E���l�Ańo!?��Ϲ]Æ�c�ۼ��P�IAc�U�1>�jSL�G�BI��E�@Ln��\vʘM�kn�E��~����1)	�$�1ߧ�UCC�;	��}���&1M�ݺ�O>OT��BTm�G��ίS�DH8�R������3F`�Ot4�p���!N��Z��ދaJ��㸴f�U]�]�7�O:xT����ij>�{0������$��՝i��#��i������s�TY��^I�c*����ҧp=Ž�a![mT熾X��R�=(����a�ø�D�?�\!�w�o�Bl��=����+S��Ol����DQ�A�"��Nw��Y��!�F@S����paH����Uդ(^WB,ɝo�^"z+�/�&'�g�!���i�x��=l�J�����b;G/�f���K�o3v��tI�t:y����;cV~�7N���7�:;bIł�Z:�iS� ��D���uyd���o�U0IF���� ��,G8�L�?wSJ�[�,K�{��,F�{ET��)O���辂���g�0�鶃�hN#�"�����u�t��P�!�r8f2Y�|ȜT��Y����Y�3쵺5�L>@φ��=������=��2��}D��}����j[��͟�@X�$�1���6X��=OAU0������!�0�=�߉H��v�N1�Y:^�{�FSs����A�2Nj\@O�*e���"= +.AzQJ����XG���˻�ݾ�6��hu�'��v��Kɲ��
p뿘6_��SRM&ԇ̀���+?���a�Bހw�a��p$��Q!2��vw��X�`E{�k����euyWü�Y$[�8o)�K%�~�\q�p)k��Q4?��م?��W�����0d��<&��㌮�J������Jԟtkޭ�W3c�ݛ�y	�E���n�-2�`��'�on�F��Z�P3��tĂ�uS��с� K6q��Ė5�0N)�|+S��^>H�4��nZlx��G¾�9��_ƞv#+�!�0ج�!S�G=� �����>��:�{f�T
�9׬�l�'�r�Ʋ���2m%�����!�a�0� �l��_4O�teB\ �[G|td6ֲ�i��&���	�|䬨L��*�$Ǝ�n%�X�ђ4���nSV��"/s�1��iO���S*v�Os%�oO��9W�F$=i~L���N�N����~B1��m6�y��fIݥ<�[٤b,�;�T�C���*gA\��V >C�l��3���T;�
����_plS74��OlI���֐?�nT���Ai�9b����r)x`��%�$������;�g��WΩ"�ʊ �S�����LmH���C�i�V��n,�=Oʦ!��>���`L5��ଭl	\xngbA:�*��x3Q!�CY(�����^ܕ��&z��N���u��gD/ȧ������7r�x�o���,ZnI�3#6
�D���.�����?�g~�Z�s�c���@�����e�q[�F�ļ
Ճ�wC��H6(��[n�K/�x�F��V��2�OR5XI�)���7Y����3TprF^xY�<r��*������xf��	]�0(�ei]�$G�Kc�R�h��i���ױ�	�H��
=su��[mV���ć [:H�a���N2�H8Ԓ�8��ov��Fʘ~Sz����꣟��Z���sJ��b���J%dc�1��_���`�ٶ��+R���T,z���U?	�v9�7U.���Ѯ�:/�GC袉�1�եr��n��.Bјi�j��� ke`39�K���z�F����!����A��u,�h2^��r3*�_�v���r���B2o.2�l�ͼ{�>�v)E_��:"��Sr�G��:������@��c��0XQ<5�l��6Fr�F�ϑ�Pt���S��׌�!�Rm%���U�$.(v���B����}QQ�k��_�b�C 6˨��W���t��F� ���L�E۫�Q/��kɢ�F|+�����UQ@�  �袨�G6��t�H��
����-�/�(:�n�D�ff�Q���lU��]���
z�*+���d3*��pR0L7�G��b�^|Sjޤ>�����L�ϓ�~���F�Y�w�	�2��!�W��W ��1�I�>֮Q��=��o۰�~Ľ(�D���kpM�a�%?�FD�Ey�,���A/��@�p���A�l&���e/h�L�[�M��n�:�VΔu;��D��Jh��e�"��j���U|���'��밗�@���6��x�]j�ڬ�2���U�"un�_w�]m��_P��>�ϐ�Z�q	ϊ!L@ڈ̖����MoCǲ����'�aR|����`d;�\R��Lfw37۫���=#��I�
�k@.Y���R\����Uԙ��)5ϑ˨#��YN���4ҧ�kB	�;���.r���K4ӧ�W�4����!6Y(�k> �ȔU[������5�o)�G���@��@��l��K]�T����|�l�&���S��ե���EP#?UH��ƅ'�h�h��+��(Yz�[��o������ы6/(G��3�����\��e�ն�Y�ܶ��Tr؀-��_���U������������xm�/{Jt(ƖJ�ƋVl�E� ?�j��t�W�G۬�OJp����t�Y���0��_@R�ʥ]��?�v�WUf�>�9}օ�v�"R�f��z���cċ;��(n�K$�8�х>I�x�I��	��`�z���X��C�V����#{CY?�@Y�S<��wp�����܈�� B�c�Z���}2��k��x�i|ҹg������5��w\qz�"�Fq�μ\��?M��d�|�:J�?��hh�-3�57�I����ֿOZpce��V�d�Iﮞp"PŻ�{��5x�r2�@C���2��-�^u�u�m@����=�[)\EȔ�K6�5z��#����O7 �U�2�p�����v��6�S΁����M>�W���:0o.ۻ>Ǭ>�쁑j��T[�c�쌧�u�v��@�����ѣM�5�Az�0�\����׽�jo�{J���m��Ӛ�}#�ӛ^���"6!n	�yzy��;��[q�S�W��#�WB�D�pC�`��8غ�bjqw�5ߝ�-h�����B�PH7W�h_��K��y�ReY�3���V�Fx/�4"���i�ϛ�qPU0}�NT��{���L3�֞5�{ԝ25~�Xe9Q|2+�p�3N��2�g���a$2�u�$A6ߒ�2�$}�ăKs��������]�4W܋�=s:=�A�O�Qg2���i��5m��mΝE��[5)^���u���}}��0�P#`/��k�I�p�5
��ݒ����t��N?�vA�\v�<��ǧ�<~�Dk�gT� ���a��� aQy����姐�r�11�:���΄��jf-�C���䭳A�)_�صPi��xUF�ӕY�#?|�:�P�^I�����sL<0a� ]��}��}�CeX�7�"3r�1�Bֿ"1�ιuZ����*�a� �ﴬӹw|����ޔua�J�i�a�����C�S��}_��Cq�i?��{�H�b/�e�A!r�+���ܝYUA������"�4��H�b�����B��M���ux����o�~Hl�������F�mR�b�5qk��$f �Y��(��l�l�^����uj���*��@�kEz����C�����	�%���l�um~%�o�)�$U-O���p:6��U���?�x`'vJ0<���/�(
���&�Q=�\��r;KGҍ�B.�����p[�K ��T2�"�	=�3kP�$�-��5�u�xk�᧜*��L���+�EQ�BO���Mn��%�(\F�!�WE�M����Q[F�K�h4wQ�� 2>a��A�x+?��̫b1$S����I/0��Z�q9��8!ϰ�\�k�{v����+�d��͹��-5S�Q
��u2�뱾gw�'��~���z����0���U�̫f�n���΅�t���.C��S���.B$��A��Z�M�r	 ��:R�b������Ϥ��#Ѽf�'�1%����^�cgy,7V#��s��is ���u�8T'5��G{+�gב��mo|�
��y䪴����:E�q����\2DMn+����@,*���I�^�%j�0�r�����ޘ��o�3��M!�=�{����/2�V�g�.oDn!7�t0�}eD���\6˲[@>���Z%Ȩ�[���{���*��IՕ�~_>���mͫ��z&z�_�a�W��Z��&���4��@F9o�-�$;�R_�?H�'��� ��D�`d.����{�쵫*�nq�ļoe������-�~��Y�8�:�n�^��nq@H�J� �L�A��<l�h���!��![-X��'�c�Y���	Gw�~D���%]ָ����Z�kO�tgmS�0����{��2�VWg83~6|���	��NrM�B�U�����c:&�G�
L��$��
6�,�2V���j�W��'���0]FhW���^���A��
�<���� 밗�^�J� �r���L����m��ϲ�ϯ0#���<U��� �h���ZB�D��mZ%A�`��b�5{ҥ%m)��@�e���>��	�D�v�����fH-wg�>mu�p�I0}p]F�8�1*_��1&F�(���(�5_ef��e�NY
{.?㹴�D��	��O`�a�
�}���`�<�Q���D������Bx�Cy�u䤙�)*�U 0ki�_�&��e�	�����gw��1#i(���tO�"z��%.Rvݟ�!��W��Z��h�z�G�ݗ����2�͸�O�Eô?=�?m�.a	8�{����pO"͹��n�>N���8 �YK���ZI�r23��,�e���%�Rb�
)��mJ�]r!�H�Rř��'�Z�1<o=�rz���[�,�~��p��M��/��z[sPrH��nL�8�8��ܪA�M�P����ۭ'*<Z��W��*��ǃ@a��4�����J%��2��$�X4m�4�����+J2�̄�6DB��I��ca��Y�_.t�d���Vjw�1��V2^JS%�R�����;�n���-S�3z|*TIr�w0�\�
�	��PQ�zFӡo�S�t�t^_ � bD�ibw�H��m/���dʹ p�ׇ<[3�9z������	���*b2wh�	lF���K�"C >fx�F����6�&U���l�TLW�do�3N�A����yB^%�վZ��b�dhP}�r��Cq^Y�B�.>~��;��'��D��p]9�FG�s_�_�*�NU���u�4#�+���N�,��G�������]��B&���
P���-�C�J[
^�8�a�he���x�%��l�u�D}�A)�v,��`a�����e2kSU�l֝`�1E'��@SN呋�|g:�^t쒛�}}0qo#�&	W,����@�g�\G��b�3T��
op����S\� c2:��`T]V�=�斃q��S�!訔J����wTM����Y�_@.9���б�s��ߪ�3�����%tCH�RF�6hn��@x���SIYx�_m
A�Iym�I$5���;�ã��:�؈��J�/�e�Ǡ���و�
v%|����&�)���Q��"4��̽���S�[���Z@'����H��.�����vh	�@�]Ј��rT!��<;W�m%�����S��b���_�q��('S�/;��"K�WkDM[,�����A0�Ό�|Y���-��������G�܀X� �v߼gߙ�}�I��n
|��ʦ̽x�T#][\u8��_t�PGY<�9=m��2�E���H�(�<��+^wTbR�c�>��	��$��J>캳l�����p���Ԃ�j h1S��sѴd�%G�hL�vW��&7��\�Y�����"
S����Z� H{��+������\8ma��sQ6~�	0����Ke��^���X�	�@�]j�1E{)���z����FB����B�&��N��N3�)�u��}�v����$o������}ǟ<
D��[��_j{G���;"�Tݚe�)ޠ�����7m��3����Xv��`q������*Xu ������WJr��*�z���h�c���Qm�g)���O��C�=,,��(5<%U�����K��b4l?�[�X��M���Γԅ�'�޼l���	W�Ng��P�[c�U)�wbK�e[���R�2�?:� �� ��ڜ�a�;-��W���`��q<�t��ǜ�Ĩ8����a�r[3�Lͫ���٩�;�kgh�����Tr �%�mV���C6��b��Kׯ���w�}˳P+�z����tj���q$JO�^��MM�d9�tz�$|�|<-�+�����K&^�c��J.��XjDCR�Wt"P���Ȑ�][LZaI����	9��~���ŹͿ����d,�ܧ^���F�2�.c�oٿCW]۱�R֡_��Lr��wX���~�t�$�:���*��<J��
c 3��]� {u>7��WBu+0+IqP?S�!;+uT��؃�+�����"��4����?��;��SH-�>m�����
\��f�v;|1s樲��4�#6s�	%c�-�k>�R��ah�t�a��@�¸�ڜ�N�!���@��6�z���~HuB���9Ƈ�V�v4��	���&�!bDJ����|Z��cQ2_=��Xq=�e���4}���tbnpFaL��m����=�L��SD��V}��2L��B��o�LS��{H��L�nVjy���f���.B�����5��AL������<����<�͗!@�39	֧��љ�YO��D�ϝ��.3#u=	�8��I���:ga�dM!%����o�9�Ӗɦ���mi�-�g�j�8zV����դ��22�py�ҥ"�[�_�V&mD���\�_�:͕�;�Y�؅�ـ�7J �>��"����)0m8�t�D�9�]HN��{���	4X�c�-Ԍ� �����m���1~� ����J�����S�W��IBd���e�A�s��.�3��}�(=�����Ǒ��"�K��F3�>�j�c~	�~�TK����\�߲��a�����:.i��~sR�S/�\��$V`�B��g?�?�@���⬆�2)�NN%�q���#1;�!���?���#35q�:�#&�շ�8շ��G�DJU@�oO�T}�i�����y�\�:;����4���C)�㥳2Z8��#��^�QX�/�t�%����w�!�)��3m*�]����5H<���T�;��r�\jE�[!�S@@�>�RP�f@��2۴`���|&@�,,���-���ƋY�/r ���qm�!X��E�rNCi$2}o���}%:X���c����(��m/���k�2h��|�q,������K�6)�w�z��ÂKV6�w��Fٺ�NY�y���Ё����D+҆��C���s���!SO�nBu���
H�C�`Nm:�$��R��=)���i�
Z��y>�h��S8pkc���Zz��wr���)VKz�{֪��:S�D]�Ӝ"�F�l�>n�� ���J����P�=A�sG�$�(3��!�joB��a��K�'�]F��<e$%��u�f�:�d[[Rh;g�����=�[��QE�ݎ\�Y}0}�9�f������kA]E	z��q�����NJ��P�(�i���Bh�� �l���NyT���l��o����$o* �	+���N��O�`�H�k��/���@8��W�R��C�����&�t�2y|i���x��8�#z��ؼ迦�f��}v�rB���7�f�������6k�/eu��͑m�:eĞ^�TFv�Z���͸1���_�ü�%�#��e\�:O0�n�2��`P���s�݄~'�7E0<z�c�Tg��Cu��U 4}�8
>\�i����muv��"��YrBI��W
��$u���iN9WJF֫!��!#bX���t��K����&�q��̧�Ge���y��i�E��V�]X�M��y��H�H���B�f8\�56�ʝ��s0���j�L�D+��f)�@���9_=p��StP.��~����1S�`ξ�k�&����c�+x�?c@5�j��D�ʈ���ru�k�Fop�
qW{|8H��T��%:�c��ł)�7:;3#���!w���Uɳq%�uo�U<�CmHK-9a�A�G��"� V���.�h��#��m�T%��ϛ�>���:܍ĭL�N���0��,��0O(�#t'FϬ�s��Q�?��I��Op�ք�>������������O���
��uQ
s����輻x�|��~��7	�؀��>-2���R�K޼<7���*���=H���.���@n�l�ɼ��q�!䁖Qs�[����%c�~��ʀ86!qC�ɰ�T��N"�ʯ&mʉ�*��O����Ao��yb-����H'e[�D��\x�������Vp���9��3|�b*b������fȹ0���͊�>�XC�bR(���M
����3�q�%ڑ%lM��yq�^�o�����P'�~���μx�X+��WTA�%+�V�z�����]�Ͼ�`9`ga�ar@��L����߽J��\�~���aQpP�Յ7�W����f[�Uj�Ę	v�'k`]��w_fr�Q[�N=�b�-NC־bL�/��Б68�g�LF	4�J<� @���	:��U�h�h����.=����ZG�r���7i%\�H�+Źӑף��T�Oe"����V^PC�B�_�+WæV,9��S��T"�Ф��5�T��ڥ�;��I�eҽL*Ȧ�\0;�FoN]Q%�O�~���z�X�r�,m;I4��,�.�s��h�놟�ݡ��ϖ�\������fm��B�N���dO��gׂJM��$�gϐ������ޟ,,N��]�c���ϓܺ��u��,2
^�4WPt���3>�з�r�h@'�a�z���W�9���0���K��٫�X�$ \���i�Eq9�'��z�t�z�d��E�b���g!��s�Fpa�ec]>������}�%h��i��m�'��)�n?D�MC�E��.�Dk)�ǈ0��X��"P�>lK�M�f�]��d�K�0u寜����n�a��j���Uo�W�A���\�2Q���w]y�{^UBtƠ��:��+��ar�����Rg�r��*u��s���ƳHvƣ�����Rh�䫜[h�~�1����?V�I5�tEt"�1���U��=d	����=�;~�-�>G!�+��Zo>�{tg���}��y�f�Se������.��Ћ۹���xSR�;���� O��_�c�;�4|ty�>ls-�U��.Z�i�$J��sv�����9���m��c�0���^�J�6��|�֖+�Fu��2���;vk�k��y���E�E�ˉ
�#m~r;���)���MGJi)���D�p�j:<�ț�c}P�b�>ԕf����'���� +��~9���/�
U��Mxn�Е�H�̳�b�<���@f�#��,q��A(�C;p,�s��}W�AAo)A�p�HU��6��O����.f*�h���>g���j�zQ���R�>qPp1�
jYt��- �vI�K���~��{�F�R��$�MJ��5���u�0c'�]��jK����Y��X?N���r����]9�j_Q>r�z/��:��	W��o�E�����*��慘�� ��=5��ⓁZ4-��	�	�L���_D(�����)DF����Hނeϵ;�R�R.��B�'a����:W1%��ˑ:v�E�F�{K{X�iеU�J�Cd8t�a�w}������[�j��x:�d>�Di��g3!�	c����cn��x���\�d�:A9\��E�-�5P,z�a��v��B4N�k;Ēb��s).$�����l�DPg�2c^
���L1�n��g��������ME�%,4��L��lD C)�� ��^�������Z?`��"lڅQ볜j�YiE:~��H� ��?k^�JK��[wCd�MOf�4�黊� 7���c]���yNGûF�xF��*t@
R:���e���ȣ<K. �],���I_�5m[q����U~�%�q�����'�I/ʓ9����	��r���KIݾ��Dl�r�2��E
�2��N'}"�!�3��?L��3�2��j�\�Q ́�>=��Zͥ�,ͥ�L)��(�6R�r���W?n8��8��H�\�᳖�	wk�|�0��#��C��ϓ������s/�*J|#��'�2P������=)b,�	B.�d�j�t�F�K��$��Qk��X҈�w$�p���Y�<��y����%G|�8Ѭ��Xcw&���@�6Tm!
��z�y��n���Ĺ ��«/�ϭw�֎����.Qmu�^-�l��ꄏ���g)in5x=�eeq�\����mmm�N~L�X�!�����cE���g��b�" �ΚS�
��*�S�y/�5���ϙJ����&�8�3��fٗ�v_�(��*뎇ǈ.\ɖ�`����X��!�}�@�b��"1�1���q���x7���6ş'�ݺ���c�
�p�Oל+���paA;e$&a�`�V�ɨ�5�q?�B�'��}m�0#�]�o`��˳�ΦdH��g��:3L�2���L+��[��&��Z�"�j&��@�:Қ�֒��Q�A�n2fw�ل���ź��A�$Yaؖ��9A�L�6	1DF�Prs �aw@�ځz� �C��Ce�h�E��F�R�K�G�&n���,k���m��?;jm�_ԮR|^��V��՚��i�� ���"� �,���\-���UGUB0��F�q �7-�9�m���d=�<�0�a����0&�ю����6xSf�);��3`D��{]u�p����"���G�P��H���f���*ᬭ�JG1��8m�$�� ��97��Ň�b�:�* 6x��ɤFsI�yʼ�1�A<ȣAg%CΗiȵQ�3�v���PEi����@����
j���ͷWh	��J�O����V\('��n0�9R�X���[���3-=S&5����3�{U����P�s�!,̧6���zf
 V0W���A�e�`�X�~c��FIթ-��C]�f���W�գu�]|��笪ךh�?��Sl�`b1h��,����lK9��G�"OV�L���'&8�-�v���ئ�]	�ZU-�f�z*��Cz���*��g!V�K�'������.�ʗ7��]�f��Db��Z�Gw��#aUĿ�_"`�O���/��_�q���^��7u��u8�0���d�!3���ݽ����|���������s/��0�r�P��:$�_T�8/C������H�?�P�j&�ڊ��`���8��o��'	���L��@T�~	! ]LhAe�����r3ӈ�\~|M���""5��%
v�)C���B��`Z^��1�O�Sa��o��4�E��|}|�1M;�N��|`_y%��9k.�����2�݇p"LVC}۽Fڵ���d�ҁ|M��H���/�fG�+ρ�b �$��Z�}z�Ǟ����~�����A��LY|�0��9�����Xvς���DF#�^�N�]	������U��������m�
q�.��C�P𶿵���~L�A��Ps�W�`��	ʲ��T�;ѸL�`�A�7��'��t��RqԤ)lwH����^�^��٭��V��/�p�-�+Q`v���w'��B��Y�z�\��I��:���	Q5)dgn��E�bѭOb3$��������_8{���~��ΞN�\l�f��3�a�"jtE�sv�+o+���Y*_����$5lt���<m���R��m��ę����edU��	�a�3����?`6?1��e���2�5S�Z?3xscx��_�je����RC�f�|`�N����u�P��'.DH�i иp�#ם����G;w�	h'�Sq(�Z��]t�!d��S$!&ʓ,jcnC��c����mk08�;[�NOy*���&��Řl��ɸ/�L]��F�Vr�(����)z�2��(v��h3���j�Zث�+��i���_�LĨ�r�W�K6��B��:����R	�Ojm]�No�[�ʂT�A������ե�q���o)s���M��Dʘ8����]O��S�:�
��V^mAH�w	��;���gu���N5[�����"m�	J$6���%��b��lj
:8S�*Y%d�KEX��1���*�W��~�]rdsq乯^�y7�v�ԫ��r�k�*��a���H�A��Q7�l�,�%<���vY��Ԩ�1@�oT�ڸlޜ���|���|�ˣ�2Y�O�H���#\mh�<B���V/�+t�Z��#��vʍL6����H[�|[Q � ���nL�Lŀ�L�����HEkd���N�SÈ��	���� ���>�a%0���ٹ��P�RT���o��

���=/�L����
�0/vΈk�t�zFգW��p��5�8w�XpeqFt�v$Q�b��PDOc������5�N��c;�#y�@aX�̭7�>=]ʘt.IUIi���L��e�un�?��:�p���z�]�>�-\u�R����#���2IO����{�0�WH���l;��CT�a!�{-W2���	��E��$��|&#��J���h�2���p�C/�7��"K�W��St��'d��|�Z��N����{��!�e�_&�'����/��~�B�q�n[f+;V�ɴyΌ~q�� �*���
s+�l�۰�}xF��|���v�d�=�j��"�-��}�	�0͏����I&��TH��)���r���r�at���C��fg�������W��3��P�Jl�1�*���aCfQ_�?��;wh�Yа"#q�^ ���d>g[�ݝ;��t�Ef�E/!�7�t.Dd������
�e�(��Q�@K�dh�-�Z�l�~t�+�%�Į��y�5#ͯp�Z�������am�ɮ��Vݓ�2�Pfӕe"ٔ}����.l5��t�R�ߨ�W�xZk�7�g�(��:aW�	�]��m��h
�"�?X�qc ���ވ���vm�� O�M�pYs9kp��e�!�T5�~��t?��B+�j���ԑ�kG����,��� �)��k���C��9��Iqp�������{N>J+��G~/L�b���I� +]3E
2��B��� M�Cm��1"��(Ղ��[����	t��Ƥ�3Xx������¼H	zbT��8���8���U���YI?US{��P�H'6�݆8�*_�/ZF^�0���������ĸX��g����^̚���M~���yT$]��J�!.
Y6Ǵ�$A���ܘ�tZs#�,o��ސ2P��A�444g�?o��2���`��a�����ݓ�nu)�J}��m ���2uT�������&�Jm*����n��'	|����.�"��L��$*�tك6_����"�"6�	�tchvXx@$K��qu��`�K��Φh���8]���$��_�Fe�B�}�'|l���$�J����Ģ��9���S2�h]�"��n0�ܞϿxY3�Q����Pu7�,\"�Y}�� Mϑj���G/���.YE^.�Z����>���i&�&a��/�y���n3i	�h��&K%cDm�@��ߺH�I�mƇ�z�z|1�;3�&59.�,5�-��Ax�H�̚��uE
>xتre4�8��g.,�2P�Uj+����0�����~�Z-� �a��1���7�J�- �S��t���r>�IT���ۛ4o��e:��S��&t�V.�������S��?����\4��a�@5�g[.� [~���M~F�."FWg�Z{����:<�KY󀉎��Zjy���~��;�Z{��m��W���-��jQǢ²&�ӊ������S+����*ZG����a,���7�	����C�Uه6$�������YP���ϗa+sB��[oNT�δ�i۞��X�M���F��TP���ON��%Y:R=�?��# �qf*G`X�:��J��"����;e�A��D���3p��V)�R�Jֈ+�;��
���:G�~2K-Gh���$Gb_g������-˵�ǳW��+��a�V� �}��Zjc� ���yzki��訾���%l6!��M)4�����?;K4W���*����vX�g�.�ۅFy
������f��"�Cf'�@�������͠�isvH��QO��пH���iEԍ�߳�N�������Tvih<���Szi�a�l�)�s�ȱ-9ߤcۺH^�֪SC����3ϳ�m�#�S�(�V���=l?��5�L��~���k�W�BX d�o�Zd��cĥ5D6^US9|�9��cM���2^X�흾�
6�@�μ����~�P�_�5��T�i��E�����!:d��,��y@ū� Q/�ihڦڞ��E��S�HW7\ /)ɈE�"���[BI�puuf�Ӹ�1y��Ү�+�t���A�9�F�Q�
���{
C��:����pCZ���z/dh��f�	�������{�л����n}��qIL��w�pa��J{~Mt
��MO_��VX
2���n��
[��~�s8]��lm#��ؐ����U�`�p�,�#ĵ׫�7�K�Zo�v�p]��C���z��,�+�i�Ŵ���P ��6�E���&��u�:����}��C�F6F�yu9�'�ǜ�3OkY��B�R�t�E�c��X�?�SB�*�����30db��-!Y�a)[<�%^��c�x����-��C~�F��%�j�G�N܋�\E���:l��d�O��6C������QD"��ս�b�� �8�n�g��&g	�Ǹ��\�ù�M�b'�7k���������Y�Ay��e�_�����~7*:+���FPj���H@���E�Q͒�=d ��^��!�?8]��p�ie�y��謷���}|̖��bv�I�zwV�H7��۔����6^ǒ-�F���o�Y|����&�;�����J���/��b͍��C}�Nt���郶Y�L��%��TT�yf3�z��;������g9'��WV��$��6MU��o+�#�ƈ�λ����F?����N�����Z���|Мi�Y0����9�O-�hষ�
v����y��Tit�eP�QJy�%O��a���c`@b����
Y�'�:�-��K+j}��'�V�)�h0�j2C�l�p����S�f�a���?�҄wD*��v���]+)��+4Ra8�3g�y���8<+���iN7̷�c�J���l��p2���8z�m֪����V����3I����r��@(�s��������(�F�8 �f���#.�`4y�t]�2�}�J|h7#���� |nɩ� ��md�Ŵ�����!����q�u�SH�4(#AQO����W�`�Yum��N�V���7^�΂�C��c�.�8<�4�;�HM[
�"�M�����C{�AKy�j#˞ǔ ���t--�5��x��e/T��;��#�^#�1��W�|��78e�Z!+=h%K1�?����Q�.2`bك�Ca[�;>?-Aҿk���8��-'�n���|����Y�Ms$%��X�?���Ϡ�{����/;�k�^u8-�]� S	*:��S��s8�.�"����{F�ĮU9I����րv�'�Ex�X�����cr��E,n�H���f�b��]/��d�����d+�MYE(\Ţ���V����cz�\KI����i�3$��-��;1xdX%4�Vʌ�����k¤C%ĳ��;�;��u֞�X@s
�L�f6����T>��?9�0@@Ëo��i��c��K*�y�3K��>��oۃ��b��=�^���G�~�Hd�lz���6}������Ŕ�a�M�?� �,_��/�3!���*��0gɱB+��,��[NJ�]VFY&����G#U�q#�B�cBT7��@/����Z�����
�@��gw�{��'ng�0L�ɟ�V�{������>�3��v�i4�F ���lօt��ND
LM��-
PgW[>rMܜ i\�:�+��n�'�<��)��'��C=��}i���'v��"�ߜ���i��I�Y�ʞ��x�6��{d>J�$tZ��n��?��v���N9f0ېކ~R��#Azi(��ÛV�z��e�M��R%2�e�?�9F�5+a�~J�4�p������{'B�H�)����?ȃxP���n笤$�}n��!e���G�vVqR����{m�%W���{�e���͕	(���/�I'�f'��i�W��F�TÖr�7�N�;��S�nVg�
��Q����Д�@5R�'M��ZI!yu�d�3��jB4�@�,<�I�G~����ψ�e��'���8Ӈ��@�pxl"�>dO�
�L���Y�M�C~⡲�0ǫI&�˻�7�A��n�)jx��?MW0m�F>"��LK|Ԃ�.*'O"Ky*����Ï��H��p�.�P��@�t�˝��R�hqv��3�4\����w}���SŴ�*�A�\���P����+%�!�u��^u��򵯁������͙{�N�M��^�Km����t[�����a��G�����,���܃D�aE� +�ꔻ35�H٨����[�N�y!어t�,f��<�.S����쪢KU��վ��[�Ui_M�)��i�fJ�[M`�4c��,S�qآGB��l�#�|�hf5�޳�	҉p���밯��,C;�-}���O���ۄ����:`XR
�c)G��A(hť^����D=וL&��؞��h�Xŉ��S��y���ȏǋ��s��*�U���H��w�FNk:���	�s�
�c1����@Ϫu���F���+Í|&������Y��Q��8}�xnA�C�N	N8wGr��~��692֓�
U:*���D�t�+{VZ�p�{�J	k��t��=����G1cf�a����=�/�s	��z�$�=�PP�V/	��$hs��>?������v]l���J<#u�ԧ� &�]SI�_��o<\*���cg<��/�s�Q�,��Y2���s���B(�+���T��2�5�6�T����\]�];k�`�r������^���6'o ��>f,q��0@��"����"hae�l�t�ũ|$pb��zaM6/��dplZ��Bwϱ��Hլq�&G��ۂ>q��f�<�$�ا�|&�oqs���bHp�5,��@תK�wPMU|�Nln�#?a���[�} n��}���7��í+:7_�(R�>�|;Ri������ژ5.�Cc?O|M�e�(|~�4
˥��Ɩ�6S�.�B��G�F͔k�
���7^J8���Cp��K1�A�E�,�J���u�
԰}?���9���AC�!�B��ݑ�[C�q#Tp��gr׌�y�x�x4�_�:�l�Wd�i�a��е**L疸5I-X;���� �|�������R7'�Rgr����,R'��� q�^�"[Y᳗W<�D�3h)�b���7�c�n�� �B�_���@��XQ���;U� <�"�5߇&�a����ſ�W+�T1�@�ʋ�u�%�r�MreTۤZ�����[�)Ѩ��wy`ϔ�*X��'�߭�\W�&p�����3��lZVA�ǻ�uǑ�@�L�!2������fਈdm�.���
�{��.T\D����E��x��t��Bһf�b+�I��Eȩ���e9����A�5�]���y��!Zn�4�����ǁ�l�;�D��Y���T6�^A�I	v�۟�O�v}��.�c�h�:����ɤ;#;�&Θ�N��	���v�
�j3F'�3�җ[X�	�Nr!�B�.�����hZhc���)����}�C�k*�2~��N��&�b�� D�#�Cs�0�s��!�/u�H�D;�j��o�Sv���F���2�FTw:�5�1�����-�Tz�{�*X�$ʳ��z̺FM�QTY�'����4��"B>�Rl�nfX�s��K�^�<nz�z����L�%"d�޶��]��������l̖�-ɱ�TM�&���@4?v�L�t�l�H2	(���1+�U�������w����W�����QB��Y`~;�����͖��S�'@��?%�bڊ Kzv���\+�)_�h�A�L���u�h�֍?��Y�s��	��Ajݺ�v�p=QHC&�U���.$'�� bn��;/;V`�Dɲ��xV�'��m���G�= ��>e��	ā��aٻ��7�0+6$�����2��_���P�O<g��Y��Oo�Oh��P��j�w�_KX6V�c�4���q&˃e,�z��"��S���Uzr��#Hr�J�X^�Uk��J2ߚ��cJ��F��r�$����9�����ݤ��a�,ռ#��Y��u]�֠�_�:�h��5�[b�c⑍�T�w��P��ʌ ���<�~�\�6�R�{4�dV�-��C���Ĺ��;�3>]y �>2�����l9[����Q0UpWs���yA�B�,���r܀?N��E�޳�������Pdz�Ų2�9�6e�!���/+��3gh5
������_0�w���d5?�29��d���l����Wxs��u��c�	�V)��\[`�r� �&'��T�>����L�Sމ8�%�󮼴^�P5@l�_�	�B��d����C�O::�X��|����BḠ�Kz�A����%���an��|�RW�3
r�a[^DJ���K���Or�����\�4�s�aY��u�U�C5&
sݞ���2t���<�}a}ڟHRw�S_~&�J'��S���<�G�\�Bf���A9Z����Ӛw�#T��$/W��+?�Փ_VE�)��8�Np#cG���y��~���2p�s��b�����L˃1�/7��d�.���{]�+�E4�ν �I��A{j�v��3
�"�>5�+{P�ז�����H�%!�ы.�]�z.0��˦�,�m~m8�'���ĥ@tO����4Ӵ��[���FL�*f��Dѐ?l��c6��ؒ�i �QjI]n�ϵq�x�
�HB�hﰡ|p���O���`��K�=��Ȱ�l��s��uĉ��^m3a�R�*a6k9��m�Qv��.��K�F�d�\L�=�=|!#tÿc26�z��Sg\��J�����#߮��
��q!�Q�"��rY�Ҡ�����5֥��Z��S��5��[��2�&{��7x�j��E)�C�:$�JY���J*n�H �����T��
_�����&Q�����2�2��*�4��%��> >[~�8���p]�o��A���S^p�Ȓ��i�K@?k�5g�kFY��n~�S:V���vU���ƥ*��������v,�H]�N	�2%���Tt�a�ޔ��-��G�LÈ�P�