library verilog;
use verilog.vl_types.all;
entity lpm_device_families is
end lpm_device_families;
