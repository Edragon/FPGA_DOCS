library verilog;
use verilog.vl_types.all;
entity carry is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end carry;
