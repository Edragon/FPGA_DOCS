��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n���C/E����xK�Ҵ������ebrh3�_ڦrsL��qi6^'�u�o���V����ܬ��^����H�tx�P�D�������tr�񡇤{�6a�C��建0锟��Q�Ʉ��$�Bۓ�-,��v�� ��T�*�X���fp��IĽ����H.�אܾ���&?��)�ܳ�������V�]��|1��Y�o��
���$~��j�e'y!c��M��"%��g)n�u�ƪ�g��a��r3�mE��~-��� m ���߉��E�H�Ǿ���~R��:@P" LCL,��L7p�wzքhk�߄@�E: �ʋD�yS[Iǁ����b~���tJdEQ��I%�A���,�l�Rn>'���G�tY��T�K��Kn�R����8�@��14,Mn0ـ�8������n|� b���k���q~�u���i�DT4.�8vx9U�?;�ˑ�@^��2ם���}��C�<��W��y�8L�3���k��>��褌��ƭ���.*u!]�|�2�Ae��# BT�@��&/&��+3~�W��_�wY��|f��Y(�΀���t#ں�oD������@��gI�A�F�C��o�K�Fɥm��'���{H0�ۛ��[�:�<��)b�ms�`��}��̈� ����eX��>&
'%e1� b��C���AѮ�KI4V6�%��f������	�Wg�b�4^a�������%5��Ͷ�I^r��L�ٹr���PIXӄ�1LJE�E�4a�*�j����iʞ~����/��`�b%n�����d��묫����L�\�_�+[�g!��?�13��Wо����M����)7���0�T� ����ۖT`�!"��d�5��*h���2ڧ��rK��z�? ����=�̳�<0��Z`�(�L%�~��_hΆ�ʋMc	�zєAV
ONs����N���Vk���3 Y��2�C�V�!V�������J^�0|�!
��!��������Q��Sj��_!����9~�|?T�@=�T.�.T\uϤ47��I�P�O�i��w3,��ǭr�ʿ��y\Q�e�6��]F\	�5T}F)��g��Z*o ���ItJ�����Dm�j��D� UĴ���ȶa��!���N��31�-IS
�QO|���J�f�f ���Dou	a4j���e�[{K���9��F R���Ǒ��iJ�HFMz�����1d7J�L��I��Zճ�hH�,����9̟���������^, �'[�s�	�Q9a3 A(*��3?��G�[����I�t�Z ���ÙY�[�<N[���> �+T����b��?�78�_H��@�u������t�+�`N�b�g�=��$jr@h3{A��=ڻ���;nU�&J�ך�^�P�+��E�Du��p9���֖�H$)#+�[���ztA7�r�a��tuz�a���.?%�_/�̇&ͥj�_�f�� �ꭦ��ޫ\�h�xI�O���3��=�		&YY�l�	�e{�*����5����ʜG���+�q��	�y�G��+AW��i���o;YF$G>CE����$D��6�y��N䃢��3"����3���U���s��Nc,���A:�j�?飿a��e�A|�������-|��j^��G;�{�9�l��H��r�3��b�\�����I�vj�82�^�h/,x��jGd��}�]{���bq]ye�o���kx��!s�1щd�3W��J�o+?�M�F�s�)r�*5d���i'��v�����|� �!�r��v��C�`�wk��z��X>��C��B�gN�&���W��Ʒ@z�Z��.�M�O��.���.Ζ��ؽ��ϖ�j8F���D@���R���*
���c����z�6@ɷX[/��喽�w�Ĕ��x���4�0U2�����m/G~���4V����a�fG//yC��w�v�ɋ��$�#�2���č�M#��&k��@ v���'(UD�z$�txq2�B����	S屾��Q+������0Vٞ �ݏ������6A��TR��|��3[�STVʐA�)�3��R����~�z��`�z�mm?�Ļ9c�i�T��h�]ϼɈ��[A7n��@�D$���y�r��\,L���)q��-�sĸ�:�	�b���E�n�Z�=A���m��T���ϲ`�-����d!����GU*�H،�N�9� ���y�Oa�V9o��.5#�^ c��n�E^bF=kS1�_�C�_c~��
@;���g.������D���3N(�w�;�x&@Pq��/@��l�u]J��<N�c���47,d�]�SW;~�fD��p����:=��х	q���-��TNm����Y���l1c��`��=��N�>�M��� �	�7���&uLIÎC:���Vj
'VB�� ����(u�F��<Z�i��b�,���l�ཻ�?,=��E"R EHJ�s��P����qO�5<�pŕ����d�(����1�Ws7��	�, `�1�.�����a5��`k%s��r��J����n�??�����*=��ל���#O�L�z@
0f�E�P��2P�#H�B���>��/�o(��hu]���*�;4�J��LQ�޻��z������Ì,Al�����B�lgw�MG���!&z�^m�a��~}�w|��ǐ���Y���	MZ���Q�}G{��~�
�Wӌ��x7mu��o���>5��l������9[6<Ԫ�8���9烏pp& �~0��"Z��ې�3z,��a[풥.��:l�������>���0�����z�T�3��k~1t���:���{[��Z�������K^H�^��.�n��������<M쇦����i0ޑ�b�=qPwE�bܶ���I_�]u��b>ەM����\6~��3?=I3�*��D�@X�6�rG<�`���xkLm��6��`��h�;��`�-|L ,)]�	1I�a��'a�`���dF"��Cz�r��`?D�q�a�L �K��K��ω@��+D��[�j���m���%IrM������/
#f����I�Mj1
}�"���'b�p�ֶ��A�ٝ��V5S�Ӝ���a#3 ,j�Fcl�!�7`X�c�d^)���}
� U�䟱~�T�*�avE�!����d�f���ʰ�	T9|������x��,�\ ���,%a��G�V=�T�a�G&E��1V�`��	#Xui�˷8b����:���f�O��:`ɴ�*+��3�奰��Y]&'�����V4;L5�3�7��QaD�">�ę���k�e�s:��2�m�Q_��}��ad$8���;�~?�i�5��d�;l�Կ&�dC̩x�s�ၩ>m3��U�Nl�w/]��o��^���tN*�M�����ҥe�������>�[֯�����꧱�VķM���%gg,Z�_;��^QU�Z�g\�4�j���3x-L?nN�Rf
�x�h֓3�wR3�sM�O��|�@g�/�zv�(�o�ϒ�ri8d U�\t�������N����O�:,�4�a��]�z���%���P���E&��2#��T�"�{J�n�+�F������b�Z�Ս[g��5��������]@�#5�Ǚ���l���	����QԽ��Q�ٜA�\!�Q�<�_������1c��b�3��e͉N�1B����Д������M��d�г����O�0�[��?����ɫ���x�ig���m9w�����N�g�K��ٿПp"R�㫄`CP��(真u���� `�Mզ��0���>]k���m�&���,/�ۯ��V1��>���c�X���R&����`���r5�w"�J�~�jl�_.bc]Y�|���T�"r�ij�@Ǚ�>o'��ac�[LڈA�qŐ�sLTu�_u�)��Q��D���T(ߊI�I*5�%Я�gk�O���}G�,��0O']���OW� �-��&!c�c��v�pi��c�څ���M~ى����~�z��z��	��!�#�:���(<�֥���IrQ=z��v�K4�dL�q��Qo�Ҿ ���v�d��E
(8i��k���wmV#��MQv��tGȎ˪���c�ۻ�7���^�o$��A�v6~���5pք�5/�%��p�ϓ�}�}������"��^�Œ�,)�mU�v3����������fQ1b�����5���!�#�js�{�T�)`�m�Pj��x��sN�����A #������v�¸cϒ�'t���\�!�>'��;�����xG��Bl��(i�Nxi��i2�SaB$����<������n�����{�~�q&CT�<�f�/�hԌ�ʼ�US�	�>��T�N���ⴻ-٢���������޶���(��Ʃ뚽��doX��7k�I+�hޜɚ�n��3��igz�xH�
���K/�涩�RC��5G����WxnM�<�a��N�:�^ۺ��qS�zgR@�a�.�Y,��~%%G�3I��= W��!җ��|Z{�qi�I,PG�TI4��#��/������*�$�֭lXԗ�L��"CSՄx`kٍ��e|,q.�-��@���+7]�u"ŗ^7_Ym���.�VWY^.�hڕ���#��{]6��l�I�����(?��1�,2^�ƀ�A
�����*��ȭ-��-��쐸�hc��6����H(�S�+	����.�c�V��t�GC��`�7#}KXw����H4�%� g���@�g�k�'c8-��)�	� [D�']gy���$E��kż��t��y7#�I)����ƥ� �V�
ʲ2�ĥ�#C2�{Ay	d1q�ob�@@.��8Ai�'M|< ������x^�|]n=��H���~y�_��a���T�$�:�T��-���N�A�,�#c���e��ٚ�(�if�C\F�h$�Yخ�?ڨ�ȍ�(��O/�E~����UWP0���CM/u~!���\k4/�;��y����?��v7#�=�S7T��PIL��o
+�(zwK*'�mN�bA�Q7�rSYam�[���q��:&�6x.I���弒�DI��{F�\���<
H�ʫ%��Ѿ�����8 �\�6tc�9A�0��b���+�[|(�&��C�խ<y�=��b����ԑX����"�[Lb���F̫m)�M�PU�$�X���u���֭���$r��5����`��3�eV�,(w�Z�u|5MN�}�&2=��ō6|2+ ��Z {&�_5�E
A��xY��� E�c�f���Q&��Z�[���@/	�?��r��U���L�,.�6M4Ѧ�:��*�^z%Q�j�9_r�}$�a�}�~���`��+�
�Pz��F�*�9�Lב��)�'�u:��,�np�<���Ǧ3��̇Ή�T;^>�D��N�/�l���I *H��	�2f�u��h�!�.����AGf9�m]��ʎw���NPFU��u/�`�i���T��d_�\O�����Cj�+f}�V�Eڗ�M���|؂W�D��� �eh��Z�pn��]�����ܔ��5���䝺��ٚ��4Tb�_�Yv�D4s�?����[b�P�C
!xc��u/��J�����-�,��`sP���/V�+DDɎ�����M��P>��=cm�h�|�CXig�i"3�,])ư��%do��ؚ4Ju	�U�Ӎ�y��p˒�g�X�&z`�h���EՑ�Y	�>A�Jh�>��� �#���^{�Q�KT���(��DoRg��v0�Sǥ%�9wMb�2�:����y��w�L�'��W�����	]��L�g��C����|̆b�֧Iwo�5s�)��Eű1l���p��喨*M3�'d���_���.��鸞��4�w�yZB4XO�p����Ώ�d=�^Kf�B¡�������{ @��MwL����1���%��2�Pt[��EN��'X^�g��l/K��l��1�bٔg����$G��Ϣ�c͂j�z��>4���>����ؾ�ׅ��T��{��}��K�V� �K���b�&���{�@'e@��'5.}]��5P���d�%��ܔ�"K�W�5�+ ̑z���q�����'LEB����_��/�����������J�'�7 g�%ET�'ޮ�N�S^f��B#=N������'^K��?�>i%�� �Q�kZ�IF�#O������U�����ؔ�ҕ��(��$FSdjl�H:Bs�	��.<��� ��6���O�H����<"~A��ɰknhc]�-��C�L���	;d9����a+(~<�*e��<�?6s��_�v9?ݮGj��y��,XT��W���q�4�Q^6��= �v�j6�ގu�(�H��N(	��D^�������S�����x�GT��X5ؗJR1�h-Nc�����dk�۠e�=2�s0�w6ZE��M9�ˈ�O��VB�ˤ�VzB��*�\��/Cΰ�m��̬X녩��Ү�E�	�' 3k.7�p�֊M�������E~2�A7����e�PZ4wz�s6'���r7e�2�RϢI]����˒k��Q��B�P����l����BδX�����X87�ß�`c^/���,ѻ�w'6��K�+JRE�bX��g�21ײ>r?��,�i�*X71w�	Y�����K��˙��Vt	�C�F�����Q�� ނ�Z$S��0�ю�w5^[x=����0C�3x�i�?� U��&�!!H��~yz���� ��+V�#kT �]���S��¹%�B�ٶJ$k�	lfJf����s/~�/σn�|�XY��N��i�w�9���-]ٻ��0�aÈ� V�16�v��MZ�k�k��e8��cM(��C��9[�ִ3g T�ݷ�r=@��z��=P4�Jtt�49������;��)��T6WSb�u�9��(j�_��R夆(">\6Ѫ��VVf��5���y,��W�\���Nt;�s�t�.˪�]�_��@ivJ?���7��#���ޑm�Kq.&�5��\��7���وӰ%�ƮA�H�ޗ�4첦�M��wdJz�z�A���P�Y-�B�}������n�|(!�i������k�x�Y��<�Z��5�����$���To�A`@Ɠ�����^���ł۟FC�"�I�EsS/�����G�����vh{�%��#����> �ߕk���T���Zg��h��I� �v#���	�w)I��v?�!�C�����"�KH����2 �d|"L�1	��64�����[�N+�!�����&��%}����}+4��6P Ƹ��4.���S%N��U�9�rwWh� S�g��q'4�&�s^���+2�����{']p!�u�Ǡ0�i���MH�P��[#z`�yƺ�1��SCR�-��Ͻ��L��K�̪; ����5�e�V.(M�9v�V����7|�"�~�K���8�@O8qh(ĭF�vX�CmU3�T,����N jᑪ��gVG�����E_{d�ٱ�J�E��^�/	�1��9���跥Yov���T�a���/ʕ�XR�s[�y�2ɶ'޷hEJŶ;��X��l������t���|n�Z>�N��~@�mN�T�Rcq����¿�|��b����p��A�N�Z�6@���rCC�W1�A�;��DӀmh��h���g��
1b��1�r0l)�`�:
i�@�a&`d���	�d���7i69+�����*�Y�q�uGNΨ�9L�KϨ=�"C��Eb��������ϗ5���&�������<|Q� ��
��0�ST-5CV���o�DO�4J�BgYb:.��/>�A��[8��[�..�q$��8#��䃼��>G�CԌ���hddx�M��K���|S~rNn���z���N�.uS3bߖ�����h������X�KH��[���?��Y*(ù�3|��b���3�Ts�9�5f���P�W��`hjq�I�>��N@�"���_� ���v,�������4E�$xHd%��f-��?�M���3[��Lf�Q	H�U�=�yE{���0E3��x�1���y#��U�(�/f�1���ї��)���I����J�⾼�̅0�}��}�����J�2� U�0����*Y��ِhp�I
�WVYas�"��@=f�gV��۬Q��ՠ�F��f�����Tx����t�ܲ�Rl���S%8e�";,��s���)�H�i^�7/qV)���*L���������S��2�NAN�����[7�_�f��5���ꎈ�7�<�Df9