��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�����[(���$��S���:L�go�� ����v0�|
5�}�9T/z\����rny��?�����t^�觅8��ȫB�;�<�����g��܍_:�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n8�o��Q �����@v?n��{t�&c���	�)td(A]�r �-g2(�^߭���<L���	RE1c���(��%�d����q�N'�XO/-lɈ0��U�b?��Z�c�������־�o$"�ԍ��ޠ~��*�\}���k2h㎬�.I@��b{�H��eL^��C{�p�g�
�����<���V���g��s4|����p�b��Y��ճG�n3l���pǽ�n�kS�sw;~lSP	q�����
�^n.N�����Tr5"�iޔ@&���P�͌]���KK�">v�B��D	����g��[\?�� zM�����9�v��=Uv������7�^�n����9��ݎt� M�H��  �K�
k�I u�Z|���%��=)�ض�)
��(�8
�;UB�@��+-�����_��T�t��7H?&Kӯ(���X5'e�b�T��g��g�
�=�[�w�Sk.O�f+� � ^=�[4�f���%�}Ty�F닣ޠflTj\��}�ǣO$�9Q����y�������u�o�fn��z��s;TQ�!A�	2��"�eB��"��.�X�0�rB�ɑ���ɠM�����Ϫg����|mh��}���;y�Mo��ZeI(��i$�l�	t	3;Ɖ;t�q
�`1�Θ*Ʀ�jQ;c
'6�]�.��@j��M f����9��DƵ��Z��5*�%j���D�V6rR��#˯]�8r7�,�w5��肥F`d�݈3Z��ėU���}t����Wq+YgjE�K L��ѕm��!����j���hD��U�!��d�V%e�����h>F���{w��	�n��^OYM�K=�:׉�2�]��Ã8�)$cX;	p	w���;SW0��Ok�{��W���%G�����:U��ޖ�2VR��<*5	R$�;�_�[�LA�_�Lr�uG�xXg�u5���+i���k�B���и�XR'��,�A��Z��ť�6���,R����h�;��4����l�qbC�õ0�e4iO���u�:�����>��XC�#m=�9C��d��!�A�ʱ�B���Zs�X �]t�Í]��O��"��zH��w��0l�\�f�']�6�poޙ���Vk>�a�$	������U�s�ε4FyN~�>�W��b�Ȁ�e�<�X�`1n!3M��F�VAդ���2��?��g��� �I�L��|E<7鏊�FV�iͨW����ޝF�E�v����[Ƀ�6��B����ʤ~�����(���yC�F�[a�_��-p�HPzRJ~�!�����|3Ϝ1a/��4�rG���*�`�x֫�V��{�က~�p�d�MB�4������6�=9&�����ч�fm]��	��1>��3�+lA^��,M�j��2>M�ZE;����dKr��L����f�%C��?K�݉O�m���$,4��nj#�g�l����9>p�Nl�:�H����|��)-��N.>)j>t}���Roĳ�7�S(��^�0pc��ϵ�)XS�`V�h�C*�$&������}>F�	_�1a��� �A��T��1Wc�mN5!ܪ(%�Hds�/�-�J�!�s.s����(;�\4�8��yP�c�8�(�
vƳ@��B����^m!����(�\���r�v׹�,�� �*�#�����N��8C$��Rhq��������$�A��$��F�~I:gPE|j�O�M E��@L�P�����
ݞM�Bx�z����6��%��E��TюF�����}|��
&�z�hT��&��"�њ��GΝݏO����%}��9G|��Q���^��i�tn4��	�V�l�;�db�ë���܂o{�W����+R�E�@�>�;u�Xv�r�7U�,��S��t"N_1��/�V�vJ���x��Z7�Y� )9uӭ"IQ��+����B�req�t�����ne�d0qZ"g�g��'�P��55�����`�ه��)@}�|�-x������*0�u�FÞq���oW,++*e29�.�J�<-P���Ɵ��(�z�5D����{��1 ӺHͿL\y��u�<I�ʊ�!-\��Q�j\sD�@}]�@�
�mP�߫�e�;y�h���_\�_y#�M�D;~m�"����s�#��ɏ�ߑ{Q4l��W��δ�a��=VT��I"ؼA��o(Wt�&��|����A,ז�M��lA�s^��U�RP0�rL�C�l'�-��0�Ԭ�I�\	[��h����R��9&|l��~4�꣸5�3���c�#j㿃��?]F	�e���[�U�ۀ�$����n\�Cp�Y�OKL��4Cj��m|����<e;������)jRWPN��h��n���x)�@�מt�LBlG�Y���]��V8:�D����?Q=�?�����!d��Z��/���0�BA����L]��;��d���;?��w��
J�^�c�k���y�l�ߐ�s-C굻��y�<�.m���3���z�2+#^�a��ۅ�~E�˼�vM<P�^��	7y�8��#N��G�)��k��=�Ϸ���o\,װ孥�QagpvZnV� $[�Cj��!�OX�u�zF�����Z��GT������$��?�z&6���y��ڹm��ۉF��b(3���3umFo>Ɖ�"5��/_?z�[�����b���\*�6�ؐ�x�8"|��"&E%+S^ݲa<m1jڽ�	Y�pw�LB��
ʫ��O��~ާ��a��[��#ŭP�-�ıE�awp/�����}���P[�U;��`��b�q��mQ3a�{��}c�d�O��ǐg�ĀdPC��|~�a	��s�Z��M�K����8���iI�1�At@T��%N�-�)��P�ч���9[�(�-��b������z':�=�Q[��/�jt���D�.�|T;����1��?]hN
=�R��P`B��:����|���W�X�1yyW��e+�}��3�����mZӏ���Ύ�{���'W�a�Lh����Rp>��R�U\�;i����>l�QF�*O������=��X��J��V2W9�7����P�%T$X��<T�q4��/�eb��W�;"/��	L��3,lZ���U��+�kt�h
��J�X���@���8h��^�x��8$7L�):;����e6�}O���\��Y��/X�J�-� 
����j�,�f<� ��ň����Y�G�0a�0�A_=#A��.��g'�����lvЁ�w>��[4��㡚�����p��L�vf$(h��P��b2uȇ	D����[�53f���9��C��g����[�:�fz�ƍ���:�E�s�n�c� X�e���9������x	`f4�7�R.)�;��x�A�OG�9��[��`HG��b	|�'�Mʿ����fmd:@�H�9R���@�dR��2wm�����f�ɞUY~lO�߽g$�Q�?9�p.��LZ]$�Y�O����N�E-�|A��)��g�tQfUY �$')�=��!�k��v�m�a� NK.�UI�Pp����>�?�1:D����<���N �l��s^X-��s 凳G*@����tfx�1f3�����Ogk�F�M���{"N�n��q%�2t��m��%�{F%�S�]T�\��)"�ڴ���ѳ%���ژ���;3�����VeQ�x��{��_�c0f|gG�}Uq��r-ս�N�q��vҧ����'5���U�ۼFGN�����m���F�C�`�C���������G�X1��?�˒發	;t�p��F_%�r�p+��)n6rR��XCN/�.>'$�
C�)�6�6h�cCǍ��,�K�}�Cx�EtX2M���,�Ƨ����q�^ �uͩ��F).w��uU��PA
�b�8R�4䆕��b�1�>���d$���ȝ�R�4k�/��=1�$�r��]I�lD��k��&���c�+#�J�wB��X�_=\9_��<�PS}�a�1���q[���t��|�::9�^hی��U��u����6���?�}�Te-QeH�_D���!q@�(
���U����󷨥)�2�q5,pK�)b����o����-����F3:؋���rI���q����&���h ur����8Ⱦb�!19�s&L�e����E��/��~�k����H>c��@�Gd!bʿ�	�[��r�J%�v�팫�ý��t�鬚�����O�(�%�����tXL^�
�/�s9� �����И��K^��a�|B:�S- %�k�>�h�|�h3������85��]�vkw	|�Ƀ�߆,+j��M{��0O�t��z��>8�nWE}����Dj���G=��,������aЊ�̧L���+�����E�g9�����Opz�-R �[Z�u�����5��1�t_T?�� �& J9�ɹޖ�1� Q���25+�>�ߪFvXp7[V�� �
<%b�{�p�itȚr�籈�j������f�O�u��Ew���[�-l��nY��̨�c+�I��Ϻ�Y-�Ubo�.�B܋oџ(�i�)��F��=�[)�Uz��R����-��� ��6T��!��%T֣dz�*�>$ב;*-d���l�}R� H������~��є�rC��]��z0p��yJ�_� � ��{W��>r��u��L�*׽�\�w��J8������U�j��3�VK���P�_��eo�$�n�b��>G�zMY���qgx��%��u���y����5�'��I��L~G�[����Q���)��=������2�#�y07)��,o� �GH#w��1%��s�v��7�Q ?���)sṠ�έ��vp��kEF�Ϡ���5:�N��;)N���%��G�b��m�1���1�]Í!!k1-�E�����#/5W�2�����9f�3@��޾�����Gr���L�Yv��H݌J�oۤ_��k����z7�素����Ŧ�;$&��P8y-r�t"qX��x�I����{�őVޅ8<�v��C[�Ǚ��OhEh7f�@�n���|5.wzӍ�r+�5�Ȫ]����S�Rh���nE��R�&N����F���#p�CN�E���/�hI��6��_�UD����-����4�m��Z��KaVؗ��ǝ�?�wAY�G��Wi��#6��80q˻�ѥ�'φ	�`X3�(�������7�����,�0�)H�{I�oܽk�a��W�I\.��sz�aFSj��{�ߑmO��j���ƃs�?��X���ʓ�X|���D��ț�Q_eQj���6�W"��n�*�#��Nԓ�N�~2Vtv_��Ft�dKk7�����вK�r�\���&�|�}��$_�s�M䌗����?��	7�~�7���J��{�GB�.�����:���G�)�!�n��ލ���8x��k�Z���B�0�ߢ�N���\��D��.P��h�x�hW�M޸��!w���o�}����V&��B��}V����k9���u��4�|��e�o�V�KxS����/	��!�n��MVFs>	�����$RyĎ9jÁ��X�������O0�c�傒4����b�%����H��+W�zS�ä��8mh���:qy�ϵr�9�" ��D�5�\��!PK�f|xM���\��6��o�TYl��T	�8B�6�c2c�W1.G ����͚�d� �}��}a��=�9ea�Q����q;���ĩ�ͮ=QC��n��^kZDP1ć����J�6r����ӁPz�5R��I�����.��ѭ�?���o񾃘�1}��5�|�Xo��C_�� r��M)B������N�>�ݫq^�G���,}�U2�sx�2�'�4��!XPsf`��O����w{�36�"�3��`�6A~ReQ��8��M*��o᫻E��~cL�����龕O�K'X��=riP��3\:�{��^�����n2b�M8�X��eo��A�;�v��4-�o�-X��<CNy�)e�~��|}��92�Z�,]�[b\'�e���䒖�� �Ɗ}���T}%RR[���{<&^ת1����2o��zںY���5��A"+~�0!�W�4��
�>��cf�K����?���;�?��֛�)I�ZJ�MM&q[v��3�ʑ�ph�S�8ABH�)�B�@2}qVP0�^�N�.���mNwt1Z1�ó+����ō��o��%:�б#��ܮ������tX��x��rj�Vsc���V����)�~Ɠۖ|Zy��T������ה�gܭ��le�a���A����_9�Z�����\��R���v��C��W֚�Ɵ3�Jw[!��'���y���P�X�9��q�uyς�k�|��VLԱl
;$('.�s�f��g�h��	�Cj�����`����-"�놮����D #`�V�bb���*��0�9��Tj�I��z�3G���9.�z�A��xVCB�����M��X?ź�o1�Kì���~��R�x��}.�4��=qoPf��c�-�<�͕A�q���	U��'��������>�3���^5�
"b]m���T�gG�$��Pxp��%u�3< H��mx����f�.7�،R��W���E��JG͸�ucA��x3�c-�,�UT�Ĩ}�!p*�ۃ�\�7��Ղ���s�"�Pn��[�"��V&��d,�V�-���$�G�ze��h�=P���	*�~�c�(�$(��0�[!�u�V�_���#�10��Ji�f]G������n�xC8/�g�B�]3a6�jf}�6��7�q(��./���EN'O��RR�֛��:c��׬]�)�SZ�"�
�A��{-�ш�:�4W��L¤J�/>A�񶽺yr���=m����Ⲿ���!?U*� ����_- �b:�mS�~���[��#,�j��2�����Uzf����9�����-��Z0��,�����~K��}H��}��Ywһ�=������x�Σ1(.vqW�=�N8UҦ�,t�U+�↏e6��m�)�������=��U$���R1s@�7S}�6�l;	��u"��:'ry%ܯ�ɳ�/��
�}���t`���TO�p�T�8��{,��ot$��ޛ�"x,&�5�6s�Ƚ�����>�,M����W3)��_P����6W<T��K32�T?�����B�8�Ȣ�N�^,���lα���L�9�\}J�?:I�ߓ�cs9��vߧ�􇂨�i%�K�b���5�QT�|���;x��!��W��⧪פ��X�� �ᅪݢ��fo\�JrӰ�Q8����We�g�݁�{����,̽�����zkQ G�b�G�א����9���&�̝�{9��T���[�� PuG����2
��D�G�|����F���-�����& _�2Wb�ӓ�^��f���U�ϲ =-�˱)�"ywG8������l����&��R@o���f(z�A��ƪiO����|��&�~�ó��t��yk0�9�nū��aT�C�F֋��1�=�������H�ɔ>�kq�{N�����L<$e���4��H<��A:�1�h����IX\�]��Z�fh�¿���	+����H��"�'F������܅��\E��o*uz�x�`��/�7Җ���_\j�[���VK��k^Z湆�����ϖ?��=�i�Da2ye�>ν����Y����8[]�Q�q'��{����xh�9u�Ť���0/*��R�a�hF(��8WB'�Q_L�́����&/1�vNX��gOj۟�t���u׸{�uSS��l�IȆ��Z����"��t3�����^�L#8CW��א��]ș�+{_)�p|`�<��H�;L�g��`$�zM��DF>y��V����f�d�Y��:N\q}�bW)�S.��A0.�+��M��!�k���XFP]���csh��;>�G�cHz3�6�.P������t-Th�-<�&x�qN �g��K�3�kE��G�v(,Ǯ���Ƌ��.�����4�;Y�u���d�!�����ҩ?-/S����$�W|b�?|Q�>3�E�>zw0�䀘e"��9��s�]���N�7@�?�&�d��I��Mv���G�q��3K�����70aQ��FUWM�E�n�U,{v����	n�������/�^��[��J���ؐ����- W�ᏽ�O_/KW�*x�t��[�dĄ�/Z��n��Ň<3����d\ΰC.�<���ܟL �9/���Q�&]*)� �c���h�l�n����	p�L��3.��S,�P�T��b�ߜ�e�+u�63/��)���&�����*sLS��&G\T�(�����H������l�o��A(��gU�_����DVj ��fW�晊{�/(/l��Es�iЭL�Y�O×��~h	�{��6f鯕�[u�ddEKȗ��	D�-��8�WtBc��3MCr�"[jO�**�d�X/\�:%r��z��s��7�_:�ړI뺉��e����C���KB�>� 姀��MV�qG&,�5Q~��L,iA��V|�$��Ćb�L�h�U5ON穰�Y���dH�����m�e��J,UZv`W�^+�d�w5�	���c��,�2�9e6�T�K�(9�jB�f~��s!���Ѕ�'������RO��������#��4I�K�P=���U��ʻ�2�<ͧ�a�?WƁ�Zz��n/`��Nì�]D��Ċ>y>��.��{���1A��5��3����vj���n5���@$�W�y��N��%]�?�[�;�Vkb��7�aܿ�	,9�j���s�P̡)�.��� ���^�>��jK��h{~�`�yd��F�E+N�h�	+�}e�
<�iY�7|�~�]Ǟz��(���q^�����#^ǫl-�����9�B�Bh���m/o�6 �/k7�)�K�VT�g��a�`E��=vP��Ɖu6��Ò���\��%G����1�/��ك�a�>.ùm�Z���u@،ֲ�1t_V�H���P4�97N=�e$�}��0-�ź܁����㸃�����e�8�us(9zC&����K�/�6���-�Bx�{�ل���'����'�['֡�_���F�wsD�n4^2a;d�SI���5�B!H��^�d�~�;BE���w]���9|�T�G�u�̏�m
�q]?F��	���6�շ�����O����J=��đ�j��h��#�&Ǻ_�������o�Z��"�z�+`n�����U�
N��~�[t�ٿ�<���M�y��8�∅�`ʅ?��o�v\Fm��Q�\v�ǲ��>և��s�� �Um�%Z[���%*y}8�0v;x��B�1��L�w�'�c<4c��僐����7�"��rm��%P�&��� I�8b�J���s٠�,��F�T���#7�$3�
�`�GC PT�o܂��]1@b�l��,J�)P^m�Q#��Y�Om�r���f^���t-���0�l��٥��\yRA�6(��>�ި��3�"�K�H�6)�8kB��&��ltg���.��~����p�q�<��+�f�j\����I&���Ђ��uT���w]Yk ��\)����>�zl�!h���z�p"3w���J��L;�aݗ7�\�#����hd�|o��`�o�. ���JX]��`�MQSD>9Ŏ��M�d��K[2���m�}�%"z����z1�����a�7�-3L�v��Fy�Jx^Ȟ��g�5����Y5�A��9JNKN�)�0����O~�"~��y��}�܏GzXw{K����Г|.�r�W��$�ס�-��c5�΅�|�����j9�$V�oi�=!w�,9Q,z���g�������{0��x�Ӊڀ`�:G8y�.n2yAϠ��sL��PՐ��X|�a�2返^��j!?Wu����`�T��Mߩ��
͚�����P�~R:��1Jx��)2-�ֶۢ����"����i/����ANO�c#b� _ޣ1��u�ȟ���W�`O������e�k-�Bk��Q��t�8�����0/̇��|3%���`���]��SG7<���/��Q���X��b&�σ��C��)�m��v��6=.�~�ջ4&wV3�Hs�]A��H@�Gj6G��8 s���Q���u�\s?�{�6�W�)n3� �w1�|H��L_��y�)�F{\P/,{�R&5T�am�وQvV�Ͼ�������bb
�ۚ��`,�q�3�e����P�N'	,�rK���u���A` ���D��뺣����ƿ������&m0�=���y�*�ɥ��_�8����^�Rȓ�����b:�=�=a/��4��q�k/i�w�2���#�!��W;̌{-ٷ��-<����y��
�]����H��Wv.��������+@D�+�N��[&o�٦�Zv����eֻ?fh7���;�$F�+J����q���+$�)�iՕSQ��{f���B�O[��v����GQ>��P4�lo�J�k�x x�xߚ;�i�2��.X(�	�WO�H��8���K���y�(����Ln%����:�>N�T�Wj���gJ�m1$�X����	�b>V\�u�MF6��D�����ǃ4�A̹m×��\5�N���Ң����ȥ�H����@�u[2����~���߻X�!�-���:�$�!�S��f�͟�?�3��G ��p�ѭ��8�����\��7�ߢ���l��U��.�L���訫�F�ETK�λ���_�7-��]��|�x}Mxn��!��`�_��4"��Lj�Z�cʾ�Bm>tF��^������E�Ǭ�Ǐ�avQK�@O3�}�x��x+e!q�K��?�k7��=��
]Iv�0�r7��c�F�����V�Z��<pҦ���`�!�`[^Z�Q�)�ڡ��U� �=�܌2U�e#
C�j��}4�H3ϋD)��>�G��FW�"�@5H��ސ�%Y��!k컿�/n�?p�zx��h� �+b���!��1���϶�d?����{�m}�����2��ԶS?ub��b�A���ɹ�FytB5�Q����y�W��,���f�̑����y鰛�GB̋�o;+�����3�`$Xq�od�$��!\�8o����宑�#�y��ڌ��Pc{�յl1�.m�� ]�K;�P<� _ķ^�����pLAg�u���'^ë]��u�o����']�"8*��I�9OC�C��1�*WE�&)vf�z*fN=ɿo��-�,i6���ĥ&0��¥㱗E�{!��e��{��L�V��LF�@V�Qh҇�3/'<5�2�@�CE۠�p�?F,8
�gqfDA������D�yAī�'>����d�{i�A�`��=18FS��{jď&��q�4,�����HK�����{i?��ُ@Q%�������>[�,e�V�K}��CC	K����a���4�_���9_��H%�tkɛ� b�!XV�y��E�P�9F*��,Z��Gi@��S&E�!��b������"q�D	zt�q�qM���ͥg��d<����i��!UQO��&�a�ӑNK�[�_Ka��7�?�E�iɏ���؈����͔C�-w@�P�Z8�`�a�Uu��Ux�a�戭��>N��m�<bge�vq�u6?���
�L����3܇W�E��j�����U�Ӊ��\���(KrRyNzMHS&X�u���"��?��h�	݄�MӃ��ÃQ�&pr�A�Q�MƑ2��$)�L���4U�/jN/ �������]�(���`YQ���@$e�h��}<M�p<��L��6�i��E�� �5
X�T�Ro��-s�43�]�:��f�$�z����4,:ߨmT�L�(�V��vT�
'�(�^�p����bӏC[kU��Z&TՓ�'��D��1���{Ņ�����k�s%���K9�v��S���1����gG�i.��hڴ���R�?��K�cUe<"*N^��Y0I�"q�=�wݸ�� 0a١�Y�5������)tP��v
R=Y^J�X��Y4*��z���U�!���b�C�=�{�鑈ѩ�n�_�X���u�8��40,�y7�%4��X�;O<P��ŏi���#$;	|n
��S��Q)�̍��Xİ�l��ةi���ݜ�̭&z���l�s�bW�1��ݿ61���8���7A��ߙ�?��C���Zv��/p�m����t>̢��+�ы��j<��Q�9��f�0$u����b�*���N�l6��?l��d���3Dn�Iw��~�V���:,P�"Ǘݨjǯ�@��~�_#�1O��+��>F����
�1#�ë
���/ħ��y�j,Ϊ�I:!}ظy��#��*+L�c`8�bC����)�Չ�8��������zJ%T��\M�w�p�"JS�]E�Ŝ,�C���G�`ykݜm�R��;�k�>z�Lr�lh�R~8�U<���ا��`�-�3-i�S���O`	��YP��F^�aА�m"8�C���P��Hkv�1W�Y�_~�m�w�M�F)Yk	�o\�#����wF��K��7���C�'w���*7( �50u���������Rwb.���!/x1�6���3u/Z5��7�\�����bi�[Aa�sYM���/o�vC(�7��B7J�x?��({� b��Ρ�{�3�����\�E7�e�?nQ��Bܹ�K����Ǝ�T�z��I8��=���g�����9�X�P�����P���`�:+0N��1�(�CǊ�����?��zb^4e2o�zI�hY��[��e�������i1�ro�sT��G����5!4<�:rֿ�U���/=q��)�)p��'�@S�íl�)-B�7mg��}&�!Ӆ�d�%�r�QR�l}é���WW�Չ�?�`�@Wg��V�����C��	�;�9�g&��9�H�̙�M���ȫJ�D�j��|�;��&��*��J��;��>:�t�w&��^����^p�چ��|�:���	d��Ŵ}u��i�?GG��aN��L��x?Sű�]��ܽQ��@�v�>�|R�on�p�N�ZG��̣iY�P�N)�?	.�����çx�Y��`(�<@� ��J�GN���#�A��s� �F��EX%$�Mr�I�8j�����t���iճ�d��v��4��F�~m+wj��Q[��0���f%����gh��T�xL��A��'I�A�>�T�y����1	�X�o�3��X���6Şmٚ��#lr�P���]e��AL�
xbH��S|�k���G'�J�ޣY��3�*9կ�Z8+� ����uQ�ل�R��$�G� ��G詴(Tz��rj�Os�S������F_b�P(�x��E��e%����v,Ξ��P�����{��!�luO�A�}��n��ƨf١7)��S�S����9+�N$x�U��/ό���%���P�\��cL��,��T�JE6Q��߈��c��T�{Zw��*v�z��zQ�XP�q��s�8�%��I�Ǘ�z@�DGD��
I�V�q8Z�̀O��K��9D�"�����:�(�����9Jw[��
� �*
ެ!D�6�p�)x��v�/vn��������ُ���c�A�D�'�,ގ�	�ȡEN�
6#�ԅ[0<���H����Cw��3�d�������,	֍��i���
��C�5{t�	�3BS;6�S6Ad�?Jg��9}�:Ģ�UhB�%
{�M���_̈P�8g�yAq�9`#k�F����_�& <���*�:/`yִ���=��&Z�f�C�ΰ�W!n��Ή�uP��2�1	9h��Ӎ'QK^�ᖒ�Ì�Y�����y�Py��G2\�K&X�i	ɟ0w��fn	��O�"[��8M�*0�2���#������ǅ��?4֛�Y��Xd�O�a�x6�.w�G��+0��{�Bpwjq[�n�� k�6}MGE�5R�=�hhj�J���}��KwuutU�؇:+퀌�ךw��+҈�y�y;�֕�Y�D�ǡ}]�xj<�b��W[�Z?m���K�<r˿ZL`����5���>�)�0�\�W�؝7v�k���\�X����fu�cx�~��|bQ���¾vTJB�	�M�/�f$'!D�~5E��J֊T��׭+�A��3�#��G����s����F����ڣB\�C%�*�ȯ�|m|�/��E4��_qK�`)޵���	_�Dt���[[ ���@��l�\��,���I
F�u�#�uc�CZ�K��3��B;KE΂�ne��5�j�~�Ԏ����&��5��玪�'AǪ^K5�>��$��V���P����"����?]n�q��P��Ή�׋(ى�<��b�``.�U :��(x��c�����@����$c�Y���Az�3C�
�s��0���ߛ�+8��w�PH	��T�t��7dG�޳��#��`YCϠH	�O�@�kj!l|�	{��QOq��RG�lv:!�P)ӊ����L�S	~�����v��O�Q�b��@i`	�����n�}A�F��|q�Q^�O5���#��f2�f5h���	�;U�LO|����I�\W�=��B0	H�Iq]�@|F�T�~����
�����W��E��Z��Ȱ��d�)�F���+/kӘ��O?Q�lH�\e�
�JE�+ܿ�5��R֛9�O��Y|����O��(��:<Ɠ,����n�I���1�ɝL]뮆�^K^��$�3WH�=A��py�j:*~��H�wW�� ��5`븻��y�5��߸2ʺ��g<�z#�+�ƈ9IB��A�Ş�N_$�1/��F@���}�>�E(@.��.�s�eU�=q����O�F%����H��`����.s-M���톛�K�A/�`��v�Y�K�:�f�kA�LԎ�����=�ڄ}H�m@�Í������{
���HF�?�(���@U��i;�K:ž?�~霝V^�h��R���:�x�̜a�Y}�r��yb��$7i���Ykf�O쫺t�챏G�U�#@{�)ܗ6��������p�Y�Γ̫��Q _ѯ�ͻ���
"5.9�2��X̓Ü�(6�1Q���!����<o���&�:�O��V��0�|�����r�q�J��e�5��p����V�U�W��8c��ZQ5�_#:�o��t�������+���ݔ�^�O���L�65S�W�e������朰~��ȿ��.?�li����%��o��b��N
�vnp��yVj��(��ݑ�'�.m���Ԙ�.�L^���`"2�AǏ�&���S96���/�/mGl��}k�L�A?B���ً�ݞi1Xi��RR�ܳlZ�&��Sb���`��Ǒ��d������{/6h�JZ��w�0i6u�.�AC!�A$�{���N�΄g�;*�vW>,�����6��!L7���
��y�R!��i�����]bjy��������������8	U�0۫���"m_�f�028�z���'�ˣ��'.��jW%�l���\�%Cu��l���B���֪��;��1�`T���+����,\���zFâ��o��~=�n��>+��د(��i����e)�.K݊�ޥ1ø�.�т������֫v���b}�
����Ø���
1��Miz�#`�"x^
.�o)?��FJ$f;J}��T��v�;rqr}N���C�y��;��U�i�e4݆�qe_Y^!�l�������)�#V��K��b�)}���"[m`F��[�f�h���B1Lhy��p�.ry�CLA���V��c��{��|��V�o�H~�y,��h-��y6-�.���
C��b'B�g
%���@�'�_����j�$Wޞ�@XJ"��p4�BjGKyع��f+|i�ܜ�ѽ�YI�(��<�H4�*I,�l"�2���=�ӭ������=Ο���\BNN,tۢ|�vsNx�*a�����]p�c?�� �Kr~0��.��Y�,�?���݂ܗ�?f�ol%���i���9�7�N���M:����Rs�W��In���|''%fvٴW;��{��_�VJ��s�.7�`qXm��n���ђ�{T��*���:�`d�i�nwY�T�g�t�p�Pm�3m5����==�;��72��Ԍ\�C�E�9]K<�,���a���F��ͪ1
�ܶ�;c���2,g��Q��]�$�z��I����]�1K��:��'ഛ����z�q����@DWf�db��UV����@��ۍ�����8�o�n٧5�'9�ʪ;c�8!*ܦ��X�@�8����SE�á*A����{�pfu@+O�7��{��#RI���H)��o��A5����!!��EJ6bN."����0�q_uq�;g�,�Hs"��g�|���ť�s�?T�𐕆�煍4�x���cE�d;���V6����ܫ�b����8[�f����	�7��@�RJ�{���M�[����s����6D�@��O�WM[}��C�+�o[|�H��B\c@���͸A�����Fj?v�˩�i�C����0��e� ?#�����Z>Ż�7�ڨ��o��jq��ad<���/ ]<�,�)iԟR��;!���a�|/�_v�x6N�wD��pPc)�����Ek��Z�#��j�G�����b E���#�Q��gH��|���V%��0^�S���&�%��Qx���&�f�����:��3yǣ�6��[�:"_րԿyE��H;^��zB�S��Bh7-39�>[�5�_���2_�)�.r�o�ȯ$Q3�����YeH�F�)��S�X
���]2+\������~�b��~"��@�1<G�)�j��r�����1�7>�����١��8~�?�|-)���)�Qv���qW��B����M��;4!���&�ȭ(�W���'�����&�p��32l�9�e�9Cf����R��|]IP��y�μ��b��b�h�@m�S�.���I�Wn��9*I�cΗ��{#y���d ��*5eou��+؜+�l&�����'J0le�V�Ճ���v�z�}��@==��O����r7noqIq
�g,�A��f'm�"fr+�}�Ϋ��:��}8(n/gY]szؔ�^���/�k��9^��i�8�[֫���X����Y�oOZ��� <�MuEX�����Mݐn������y�rz�o%^�/ִ��<�]����7�h���&2[q�� ��/�
7=-�!'��k���˥��>b� t�,���d�s#"V�"#E4�~]}�32/�թ��0���I�����ii-��qw
�����5Y��?��t�5g�e�ԻL�]���!��c�f"��ZN�X�>~G��eeKxձhF/O������l$*/;��H��AIIC��LSݯ1���Ң��'��[��9FZH\��oЙ��J� 	��f�i�~s2g-\�iM�2uk�Y���|�f�gi�@���L�)��������1S[����=o7��pY�v������Tp�2�ts����P�sx]�>}we@{���l,��ڄŊp�?��(�����轩� Kc �V�T���$�Kc�,̗U��h�� �]	-�sr�l�j;Jv��[{.��D�y\ë)�jV�y`Nv�yI�)s�.xԇ#h��*-�'��<5���o�sE�2i�DZ�	�M�YJUFd����R�M,�x��B^�'�c������I��z���؏��j��pҖ�=��+��:�>ȐSa˞�@���UY��S��i�r�}}h2�g������T������+Q7�*�씔*��v��WY,i�܃��Y��A�I�& 2yc_��G�	|�p�%�_UU�]�xx��߀I[g!⁞�$E2��v��|��з�?��3gfϵ!*9[	%���ѳ�e����#Y3l�Ej �b���	f[L+�~�?b�P���<f��"��rO�̔�;�t�y��4>�p_���	�h٧��n�1Z�_s[��ܲ|g�7�%��n�ͷ�ƃ��R�`��1=YN��ҹ&�-�=lq������.n\��!�i5"f˹���8�� K�S�q����o_�� ������T ���%� tpnN�
.
�X�ى�6~����4%�DB��5v�*�=x���C��+��Q�t�pG*�@"*���"꼅`�'��^A�&��ěU�C�r��/:O�tb���$�j�Ȁ�	|��%��P7(>�Wc2C��r��bѼ��M����՛,ٽ1�b�S��U݆�r���H��+��(3Z�ðȂ �4W��C��|�#��[�B5H�{�_s��R.��N�îP,�i 4�i]]�ї9�屢�T�?<��5��x�̑���LE����2<4�V]r�'V��gG�,�8��&X�E��>�.6�@F��;3>r{�9jB�T�2���>DRyiu�"���5��C�;��Tlb4�Eܠe�����O���DM��N�N��6@n���o��0̦e��B~��I�Kh�Z���Y:u�� l4�2>C��d?l"O�;\��.-	� V��G���u�b����,04<X��0�����9}i|1]J͈�S%N0��v���3����%i�A��^��c
�+�{zO�<����$tU�/�zޞ��-��H�#W=i���z鯛�8\�䖡�m��^w����4/̭pٺ����;9���jD}ɒE*P�+�[�$36r���ݹFH�"%�|IT�ߊkH2��\ ����Cʕ��Su�g^*x��������xV���<����,`�	{���/����  $�r(���W�A�Q{Z���׀r�/Q�� �M ve�^+Z��47LL��h��zC|UC)��.�) W�s۞����S9�,�P��]�&ec��c�ݠ��P`�>��ق�>	"9�G2��T�����⢰<��D�z�{uC�ڮ���1� 4���]L����V��i;ݎB�}�$q��683À�(a�U�g���l�97E!�g�9� �Qcu&b8Xo����+�4˹g�Q]m}6颾̑�����U��WZ��o@�E�Li�K�X��7�^��D;�h]xU�{g���Uu<����a�#��E|�*-ܝ��&k3�!� x�ڱ"+[)o�H��,?K.���_%��Xv�����$~���3�"�~��c�=.��؆�s��K=xIo�D��,�Hy�ǒlJ;o'�a�&.�������4��1$��r�io�-;�|�KGׅ���-����f��~ɩ�43�������t2{�Dן��9ޜ�㷃�{�����o��0B�(,��n�!�S�$�t�1�j�bX0=�@�c�9uԜ��EX�26�&��U�r�.5�.�3Ց����'��, #i�E&O��.�����@
�i�ֺ%n�׺�B��('��	�@T5^q�ХZ��|�����ޗڎ{���qe�	*k���@�ő����:��W�C��"��ZǄz�ؘbQ�Wľ'�֮��Ӌ����"
��h�����?��(��c��\ͽ6:峄�5З����5"�j�)���ł(am�^˒ߞ'+cRɸ��MT*���I�`N��������V�=�����i!�Y��!:B��Q�g��k�P
�8Y[
h*� �VD�/�C��v������5[�WZ���z>�?]��Z��ɮ��W�1���N\H� ;cs����ww��}e�����˅��A.������MZ��@�H��p~�k��vD7�&TM���H�'�s�5�l�A�J�eb������|Y�T`�?y:�rzԃ�O s#)6�%�d
����n��^���a�h�5nh�8:~�Tf���ls������u����V�9� ��I 