��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�����[(���$��S���:L�go�� ����v0�|
5�}�9T/z\����rny��?�����t^�觅8��ȫB�;�<�����g��܍_:�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`nq�a���FU}�a��~��;C	��ӏ�)�b�"c^ۻ��12O�r�T��ݔ��k�mڜ�øw�v�;��`��$!��t�C� ~���u�+AZ��s
�g\��F*Y��mJ�tb咣�|%��!��h������+7�v!�:���L��P��NbFB���kٜ#Y��/�S�Ay{ 
ҎP&��:�=�o��w�UAW#A�d"��'r[v!Ho$ntg�b�Ah�"_`aS�xj�v��qu^��\�X��؂hYHB��Z���%��~�k=��G��Y����A��#�4�PH�|�����c Q�hԅ+qB$��G}�j��~'Q-�3zN�@�hU��65�RU���s]�����D�c�Y�n�c9v]y����b���'�b��4��AI���	��:����z2�����f�Œ��Dh`ѐ+�L��M�eK�I�g��� �Mv�Js��{ n����3��4N2�L.OS�yOEK����H2�'�Ч�ҎX���,�m�LF.�l'�n�TYiJ�zANB��ogH9s�m ;�U����Y�%�.{Oa\�j�m٫���JT��
\��PU�x����v�B]O�+S���a[�HVX7�ͩ�(��xܘ�����޺O !�QX��j×��s�h�����h��R�	opE�᭕m�	�g$t�[�������8Qsrxf'�<����&�3O�`�� ��:����[t+���UJ��F)�I��UHts�ܝ[�Y�O����=%�/��"�ف�����
L�b�?Y����v�C�j)�*,�7Iǂ;���=ѻ�vl�c���͙��0�s�&�&��w����Z��a��D�����?�8XH���VK@|C�b�R���s٘f�;�9S��U	��<�ؚn,i��85S�y\l��O�z�\'�!�Wr���X��48�y�)�&�+�`��5EȮ�O_%����+W��C��84�8�&�E cX���bT�0������a��#��A!'?Yk6.>38�o�e���'Ə�D� d���u#h>p���X*���q��>�e����~v!�#�O�$�JyL.�7��M��M��:X���xx��e�-G�%"מ0ՅԒ>M;댊J+Ȝ�G����Ĥ>��(�Rd`�����l R�����0B�"��tܤ"�I��=4�_��"�w����Z� /�`�鹃�\-+z�-��2��{���ۯԥUQAL��UT�J��� �����^��n[�
�c��[�U*O���m�Zm��'�Hk�8 ��V�/�Mm9 �[n(���@�F��_�G��
���N_ ��a$PI�*��^	f?��>C�����:Y�*x`���@(;��J6ْ�*�X�����M�/��^]���Ĉ�b��9��x�"j̛ ��Ya���h\e,��&���%����u���v��<SU+�`p����%�'��� /H��2���gV���@-U9a�R`�Q��s�<����NR���{B�+~�/�z&ɺU}�e[�b��S�I�q���/������b_g��7��e/�s��#yt���\�����S�&#�G���a��ZAX��N����}ϔ��ߴ�Ҹ`��#H7�D�Dg�ۉ������v�� ����DeT7�I��ڴ4vi�@¥����E��ՙ���:�z	�[
�L5�	�VS KK��l��5mT2ȥg��p}�9Q�θG����-���^�翫M���D���C5Ap]�_g�s��bpE����G��\<�����D�A`䦡�L�F^�SH�@�J�#��Ӄ��� \�D��u\;a,F�/���E�.i,G���-�w!�3���\�z:\j�9�_�y���b����6(�.;7�#X�Ϻn�/��NY��Qt�����e���Pf7v�Gy"�\�ݛ�a� ;��z����0�D�bm��/�`�f��G��aF�.H��Jl��"ƽ	�-�vheZX"�H�"´3* )[��ZF��um�_s�K�Kth)�j@���ʴ�]o;��r�oɢ�W�I6߅T�\S��{�c�y9���\����Z���3Y�^	����9PvG60)o�bn�����Ֆԏ=1�+��4��l��;U~�%T�H�t.�
�{���� ����9���ۦ�w������%Z��7Z��qH7��O�ӎG=׺X�S�
�7�d�=5U ���P��3Ï���fq.AD��6�>h �����U����4����l���H�H� ^� [ �8�	���*`�Fm{%u��ց��
�v �h�|��Ƴ�>o3�ǎ-���Yڠ���h��v��6��R6o��`^L?���z	6�ײ>1����j�P�pol��whJ9&�2�����	7����cοx����ǲ�չ�R�_훍���ݤt/L�V����Cl�U;�]�!�L���!ULG�x�?���GY��Q���@�B�;$�@��}s�����9r_�츛��/m�C�?z d���l���e�Z��M�\�5�@r�o*UJ�B'�_��G�_�r_��T)pG�2k5%�tў��v�m��YU�|*L��\9��3�x	�
gK;�?u�t�-'�kT��N^ER��鴻������ŦU���%A&�	�磶fU��#�Qb��E���%�࿪(�K� ?Ћ�=�ur�Oަ 2#1S��%,15���U~�N�� �A!�W��G�~����7��%Sy'/�f�f���m>��/Ũ����&��x��<��Ф*��OV���lt�O�;���@<M?]�#G x\w��5U$�ИJ1_�*�Xc�H*#�X�N��	��&�M[��A&XnU0�3�Be'�ˣ����K[�։4lRo���
<��Ix ���J(M���ѯDU�.��#t[��5��U��9�裒F�?o�Ar�����Io���H`T�`�_H?��=���^�I�dH��@](NJ�s�qC��?g���~iB�{ ����b���B��e����`f�Mł�޹)7�r�T��zk0�i�*�@�\�U(���}�J���9�[�+3C#�	rR�.�"B���)70�Y�zJ�߶B�j�����/fqol��Џ�Vy�H:@�K�������BVc���h.YM{I��5������F�U"���E��U���|r��[�;�#�V��\GoY~�G�Z_ߙ����e��t�& �Y�s��&ai]����W�+4���:�?�;t���#!��D�Ҁ}^v!��(;�a��Ym������"F���\Yy�0�M��4��A�]Asݍ5Z��T:L�Y�䪊\�6ց�n���k�rE8�n���h�� ʤ@��U��#~�Y���"��|�}�
��f�L<�����+4���j�t�8�Ğ��P�ߠY�̙T|��M����Z�<�NAL�C��k���E��� B��[	��I������{�]�o�o'�S�x��my�^[H��S��67�u��g��C�i�lU�j%������C�lA6�Z�d8a�@�9L��]p��S	f4X]�$ł�P�$��������4��.��2�U8o��N�j�t&�\�VQ7����Mx���O�P�u��Et�u������s�?���m|{^v"=	�
=�;���]	&.j�`D���d�m��BY�@�Ԉ[�l(03����@���������&���-�,�jk�p��LȅB��[ �@�c�p<:�߬u����ϟ�<���m����Qte�����(��h���o�d~X�,js�	�.E1q:,p3ڃ-$X�3� `�� B'�AG8�m�Q~���J̺�5��]��z������r�7��\z��T����<Ƒ�"=ǎ�p���M��Knr�{�`�z*EQ���lF�%?��ʖ��)�z�¼Q�X��,كT� �]M��q����|����Le�3���Z��\���f�h}�����O1�v6��{��}��P�!el:�Q���H��d�!�{�t �!�`�qΰ�Z�1PK��kpn1��� R+�?�9b}H1� ]ܵ%�=٪� q� a8�f���t������`XM^H���/&�8"`頻�[�o������@���Y���rk5TE;�[a[K�6%m�(����Z�=��D!�0X ,��lؐ�+���"���9�� Q�8:��8o5d�K.e"b]偂87T�#�K�r���c=�2�ظ`|�H�-�DX�o�YD�
��8��Wd�M���rT�� ڙ�b`���rI�¹������(�A��_�z���LV�R,t�[�\���wlBkq��$�6\��/J�ԫ/���4=�+9�u�ݡ���Θ����OϜT@��I��i1n�����@pλT>��onT��)O��y�� z���aֹ����<��{2xZ(��$�>R@�-����D��t=h���[��/P����n��y�6��ڼG�2P�@3
���ȼ��q�X	��L�����Q:�����yZK�4��0}1.wb,�:Hbub����(�y�k��S,h��I��c	�.0a�Ñ��D T�F�Wv(���%����ǜ�s�RY�8T�D�f� �ӧ�i�'16֐Ǥ���ѻ���v�bk���K, �Y��.�δ�|�k��QXE���i;۞���4�b -�Ψ�ټj�ė'P��ڙɱ�����/2݉֌@j@���՚u���3���dc7�ht�۳��,�����o1��_�m���ob}s�ʌ΢P���=���,��7ѡ��ۨ�p-.	�5v���I+
po��H`�Q�_��K�/ ����띱Y�z��=�o���:���b�+2	����T�x�|͛��>�4��O�����+Pt����'���O�k����}�IV�{U���y�櫤�ί�D���ϻH���jTQ���MG���:]w�ev���>�YIـ�uRC
j���(%f�)����x ���ҌB�<��!�nvީUp~��v�`�jNA l^x_��ॸӲ�s��{�|j�c����\�s������	���1����/�a�c_�o�y���1"rk5�t@�&�N^I}��
ݎ4(i�3=|��5v��u=�=W���C�����Zq��6�6@�R����_��c#$gv�g��$��"��kOw�+��ю�Km���c�6�NF�\Mo��J���mo����-��w@���k[�)�a� ]qL���ٝS��z��������m#�����^�*3�'i����^)s�C�+�J{1�'�6���Պy}�?Ts|���k�s��LV��aQT�Пp�f��S^4p뙥!1
�D�b�� \��q�z�p�B��/6�;����Qc���6��K6�nj�a���	�戤
�n�5� �^��ޏ�ԭu1��\x����O��AT��=J�c �qB���W�m�[ZL�>�޵�~�ѝ�+���W�[��u]�:ǘy�)a|f50��%�7,�U���DL����߾�6��8�+�^��K��iK�5� 4�'��pH�a�+���^X��Y�8��j9��G��݅V�R��v=��Z���[�;�~7��������^��q��e�/�����	���`�]1���t_n�g9j�� j���"G7����W�5��x��k-��%�#��Z`�2���"c�G#k�S�l� ���M���\���c-�t��ߜ1� �{G"�擨�dO{��a�vz��ٙ־w�5��-qh9ؚ�>M3�DZA�Ue�YɊ�����<��O@h:�L�HD����^ݛ��S!�<h �.��!/��=�I��R�ikjP�[EcC�ZU~(��#HS.�,A}]�I�0Y�ٞ'׮�ޱT;���JvL��,8����0{ ��VU]=����L������V�ar�u	�Y�w�-�v�}l�"Bڬt����T�x��2��`~�˦'����b��'E���!9�M�s��7��tL=���l�1�����G1/J؆k��}�F%���������J�s32��Z
n��F��cG����DD{X\z�y��r���^#��s9�Y��,~����U'.�c��uizP3�_^�ӵ)��73L�lnݏ@���4"��ޕ.������+K�-����~�_?_O���z.�����"�(��^)���X;����<���p-8<�F%���(`�������W��޺	�M�d"�Q���$��%nuИ���\��CKw`�e�j,���b�)����6��,��C>��󜛻J�X��KEO5��	�zA_��=[m2ת) ��K�N7�4�<���%#��	�A��{�"�U���S�F�71��LdY3��5~��4x�-Ԅ��r�]�)�;��{aK�v]�Qՠd�P�lؘ�^ cc:R�Q�����˥9X�B�C��/ ]}K���<�쑘hU2�����1�A/z�AGۣv����?e>��0��߭�ōf��Ҟq(%:i�/yn��i��l
Qk�_G]��
+��<f�@��_�����4�'F��-.��֌�lWT	�(ac�*�`O+y����O�їVA��z'�����*��,
�2��a�gY()�'��M�1������7�����D|�)��2�ں�}myjJ0o����5�\j�t���h<a���lN�*E%P�#W���i�	Z1��8�=��R&�j�������d�!�{[tۯ�:?f��4t�.�99�N��΋�����)SD7	���'�������d�(���eO7{!���̥�BH�]�p�F�Og������\�1������D��`��uUO�Gafn6,1�K� Ar���ˆ�B�C�$5���(�o�ӈ�/�܇�n��Z�g�&�E|�J�Lc$@�\Ŗ^������\��aɚ(��4�̕���Q��n�(Ģ��[�^>�oV�L%�7H5���D���my�,BP7�	�O�/NS�c��#ݮ����7yX�s�.�o$��J���Ӻ�`��N搎A:�r��ăec/�V���TDNMBn�@.��K�D+�c:D�q�	A�S�P�1��G墙r��!>m�e�V��:璯�-�=6���R�Bx	�� ��|#��~�F��#�H��~��.��ś����������$Q<��~q���5���ENSh��'X��f����Kg���	%��Iw�z�VE�F�6�0���j�R�y!�'5ĭ��Z���BD�bIE~����wU�ha��������Ǳ~Q�8G'D�{�S6���w�C�����i)���\Br\�tQ�V)۔pA���xEʄ&�`':�x^�K�9���n ��i()S�!��H.֒�U���ޒ�c^dIt΋��	X|�H��ho�����<�-�R�����9�=c18���*��en|�=i�9Gg�j�
 =�Z(�9 �@�Bp�{�qxG��+u�v���՚DZ��7u���݃Çu�G�
3@:|�JE�TfBRmS\Q��갻&`��8��̓�e�*S@X	�4Ƒ˲-0�����4��>��r��]�	K�x߼q�)�fl��v$�?����6�8�k*,�����-o���K]&��N<�Ķ?e���};�{ 
��a%��V��ZvqMVG\�C��[��KsQJ��;��S��h?AμN�S�Z˼�C-��H�B�P����W����K��Ŵq�L�ِ,}�N�*�,�t�G�/�E�@ن�?��v	����.��_�k��0�l�w�Q'�v�|o�Zs��qxO����Ӌ֮p�������'�C ��T�K�p%����G�P�8��.����4rU���a4v�����Zwa�e��C���ɡ�{�u�_�!ӗJ����G�,��Lvw���*���`�����)**E�M��u��
��G(5�y-t�DmS��9N�Oq)��>��G�:�>6�[��?t��5��@k��-��"+3�(�1\f�롤t�U\��e�.!�c��@]�L�e9s�e�pw3�@�6;�{R�N�z(����紒�� }]���p���l5�2�f䲾�"��%}���.>0o�Ge&�1��ΠɈ���y�E�U�Vo�\�����Hܔ����M�(�(J�+-F5�Ch���ٲ�=�x*�\q>�"r��`������"=�(����:�fm`:Yr;KkN�L��V��F�Q���@���\g�:/�DG��?7�C�C$kbM*��R��痍�X��!�'�����
��: �u�0�6כE �0p���#yk��zW�N�������C�]�ɮ�!Rڱ��=�K=o�c�r�j`�Ў�g����@����O�,Ϲ��`�߽m>1,��cڃ��oݸ�����gd;,�põHC�u��)�g�Ȩ!ef�tߌ*���KW�O�?��R�-]|5SR�D�����J�Dkv	MG�1@`���p�ﮘ�F�T����(�f:�j��)�M��>�U�Aq��j�vk>O��{�z� 6x���Zv��q�S�s���t:2ۑ�	w"Y�Y�L���#CE��y���a5f5\�~��D!?�bnaXs�Ap"����d*��c�WV���#����8����q�grt��*	H*x�!3��j,����^���ux���1�Ty�W�e�.r�{��{�~�������ݒ�.���-�mZ{e��V&�ko:�4���/Z�� �l�A���.�1���Q�� PqV �燗�0�����D��@��$����Y�����5su���8����ႎJCk��hZs�EW�)gR+O��M�m�1����_��pm�uhohM�/&��/|7�ȳb�X~y��E�ƃܧ^�$D���N'�T����t{,�{���nMD �U;�44׼4������q�;>�i���c��� K�α���⵺��װM�ks�������喧�]��Q�w�r�1\&'훈������ª"d}*��P7s���U�$�vF��˛Z���:�1�)��ۿ��z�����ݩ����]I�&�M�Wz���U?Z:����D��L��u|�l>����
���U$$�C鐳��&�����//�-ڽP
ǯ4k8��� C���}�5�&ζ���0�Q�Ll��ﮍc��* e0�GX�s��i�b��m�e"z"3T�����@r/+�����C�+-����\�����;]� N�;E~��N�%B&�{l������n�H�4�J0�4���k�I-1��(�����m)����ǉ���&2Y3��y<�T&�0�
���$3�F�$�����t��3����vB�G�M9)�&э�۲dӂ�yI�1��i��=6�!�5��R�Nyi�T���!�CW�:K �w�R%-m+�����Hn솷~DR; ZĹ�Õ���6R���l[đf<Ӂ�~�olf)7��"xM����<r�}|�]	��
��i�K��������QF��@ɔ��5&�t'��f��O�@���v�y�'�^�`a`�]����Pʾl��6�MVR4��Ȍ�6��`P������3�,#"�%���yV�S�H�i�I@v�M������i�� �丸��sؑ;V\�k�Exk8(��� ���jd�����;h��n�[ ��N�u��P;�/��nqҕkŨ+���z�:  ��z�z��޻��~�����.���B0��9��E"Ye��xp"�'��j�������΀�oH3K�nȤ!}�^k���1�b0�3�58N�@3r�Ry��)���*�s����N5);,P�z�,{�f��|7�D�����E'��J��e��Y��m�����2��@(�̮�Yv@��Zh>as�r~>�����4�>d��sS�:L��Q��Lx���ں\x�d�%_B_]ܨ| �(�ְ�՗/��Y�%�b	1�Y�2|�QH�*���P%��u�(��»ov��p���r;4t-Z��'�*0@%=��η�\�u�c�O��5�w��ul��n�����P)�M���rͭ�0����ۻ-�;9��w���3�F!�s#���WėȌ�w�r�/�|_�{�=s�Ѩ��p�4.�V:+�&�q��i�[�_x������=$���Xi��G�!�X
��<_���9Mr���Ma�0��V3�p�;��2)��)	�ZP�87�A�-,m:����kݜ�v�&3��W�o'���.�(�@��I�%�� ��,>f�[-T�$�N0�%��($ WM�"�9f	�9���#!i�P.�ǧ��fE����xc[tvy��Ɓ3ΌQu�2*w����G��A���YI>�����d�֘��aR�E��@\d���Ԙ�s��w��u)EEP�Q�A6���,�;n��9�8���$_�ſ�����k�+�|و�W4����E��j���Q�a�����z��#g�U���Ǖ�8�5�7S�-t������V�	�U�NA���y�����)�3���*��#Ϸ���c���1gX��j�����߽?"���&i
�l�L���yݓ�G%3j�+4�L�p�4��4x�U���{d��/p����'~��܊io�p��;H��3�=F��5�#o ���|�N�ljL"���lA�
<G٩�k^_ZbM,��<��ܹƈ��o�K����@���@��� y��'��ǭ�K.�@�	=����<�M��n����,(��@Xg����S�awWdb��)6R��hהUeC�y�����'}�g��'��~R�%DdU�!i��O�'?� �L�����r�xBB<���?D��7W��.+�p���9��Z�{�csY��>�ߐy�!��"T��}�'3�:���!
�����0ܳo,U����\��,���W�6�G���Nx~R8�	��f��f`���S��Q��Z$T�%�	�߆#uq�H�A��m�H
aL���թ���훓��+�*�㛼��֬�nc�{��=���b���m�n�����y�4�d�LL4h �T���T�Q3K�Mu7�֬$�μ�i�w%��yI�(w��3��������ʬy19<+��T��Ԁ�^��Ɗ]F?I;��̜NRa�su�G�N>��ߨ�1�<Vq,~[�l��<j��Jw���a���t�D�L�m]��'(m��6��#Qڤ�F$H��Q����a߫d���N�#];�+�z��[���ՠOQ^b���Sc�%�,N��E��4�5޴ٕI�+���1��,�������{�5��+�hT���,���o�uG�AgT^{�#Mh��jm�(�W�cijn����2at4E���"�C6X{j��)(d&���N��9���<��V}��ﻈĥ_��N����Ǭ@�|�7��qQ�~�H��F��
O��,�e��:a�Ϯв��ت�
�ꍱǟ�w릓/� �r�����$p��ǊLА�����Բ�2�r���q�kq�ț�ۮ�@�r�r�
���D+��Oşzұ9#����৏��։<d�_���$��<����H�S�Ew�j����D��zA6{��8Tl�=R㷺E\OsV�h������q�Sa�~7'��I�~%��j|M�����V�]��ls=1��j�O6��v[���n����![����0 l����fe���+ҙ}*W���\{�&8`�>Y�G�ǌ���o��*��+��[kt�9��w�w��>���F�O\oD��Ǌ�6, .���Վv�Z#��O�~��������3��\�1��M���~g1��yc����2k�` kZ�#8�n-z����C7A��&6dǲ�u�sǷt+q9��u���Ox�c�S�_(�5ߪ���Ÿ�c �����Q�Z��T@T%B��ݟ~�'Q�$䝵�zR뛈��QE'��eA��g��{gD����G��dW��]�{@�a�`�m�t'�$�W�e A�';;��/5�"Y�9�|���&s5�[)u
�RP�ʐޝ��t�L-���Z�,󐝴�U���[����r��(���}�AL$�٨'w��Sy����
~Cdx9ރ4r�w%hJ�RA^z��(c}\I���(�mw��vp��e��`J~."b#���N���c���&VI��/�{R��|�Xm��\'�y��$෧�}���&�5�u�$���KOO!a<N˰����:"�84P�ע��P`��b��ֽ��];b:����X�Ea��?�z���EmpD��4��ޙiX�:�<��KN��'��'mp�⚠���(��E5�{��=���ҵW8:Ee�9����8abW܍�n]��4��c�ڱt�I�4�7c˞���Bqo�	�Ӗ���u����GW�4�ݧ&�=	y�W'[����w�#�"GsO�Hjlg8K����4:�_���Ҡ�D{�y�����<$@"�h(�<i�/£ڷ<@��c�c�[���"P�Y�"0�z�oL�z�t�G7��+ga[M��҆+��}��Q���1Q+���%�0��[ӵ�Ӧ`�-^N��E�����z��� �<�!M�k��?*�#4�<���O^����sH/&�ۨ&�4�s?���5E]��X{'�����AN@��M�+�;cr_����
`����2�{��,� .ަ��6�v����]O�{�;�8x5]�)�ً��x���a���@pȝ<6k�#?�<s�>b@�;._��?��<l�5F+�D���jd�AZ��l������;�0���Ԝ�I��>%�}��H<� Vz��JB�`�#��5j�����La�:�Kt��Q��w��9.�e�ܽ�-ĸM]!=��gj��/�V?X���Z��9g�%Y�Ǟ��i��ٲ�yѩ�%��c��ڌǿ�$p.�AO�����tg�{��&E&᜹ti������ѿk;6�*HܝsP�P��(�"���}E K�+c��8���M���kbo�E��ȯ�"�!
c?0)~�:���#���,��k�w�d��	[J�������@�&�uC)�+�=�_j�]�*+>7����i����6�a���N���,�p�ԅ}�j2ޏ���a��9�D�OnSő1,�@��TF�Ԑ����UB����^i�\!}������\�	D�5q�BbCy\�ƹ��B�������|�3�4��Gȧ�g�U!�co�;+��܏v���D�0o�ҽ�f-o�y���A���г�9|�j�55�sAKse:��/5��&����O��٢fGV�#�I�h�����>�s�Vm�T�9*ԇ�:�ƅt�v:F�5!;o䒶��w9fM�BRp5�J�6IYa ���C���II�z,��犠г�P������@��'�<��T	H�cqMO/�4��יd9 8���/P�y��^�Z�����J�qʵ<,��9��-i�5�ǦH|�n|lLe�QȾ�X�݄l�� n��/�^��53�v��G���RF�UYo`#���G�n2���:&"�wl�W9)&��%tS�>g=�O�Lړd|���ŏ#ܓ��%�v�M�>J�K ӡ#�v����y{���1�s�d~�#�RE �D��y�}��+�m>o}�$	�,_~]����LD����B�	Q
�
5Z��eeB�`�d��w���*!�g���@��=�}5�,%5���Y�1��ԫ� 2��O�N$5e���^3�F��6+F`�̰�.D4��z�Z���˕�������3�z�O���/����j���Q|W�ؗzƨE2�i��x���G��տ�Gm(��ޭ����]�
~(�_��W�;���R(�7��+���N^xEó��!��<� `�����v��W��%�4�ٗ�?a��	3D�Z��<�D
��sz� j���y�����Hd���c��["�M���e��S��ѥ���G����E�Z<���V^a~�����bC	�v�u�<?9w!:� 7�<Y!������=	� ���r���Ćm�F�&�I4��q�/�z8,jCh�e�v�tw��V�O��Uh[�+K��T��?M��C�]$P�z��i�	��	�	ϩc���V ���Se�|�xT�͙�D{-5�c���ev��"JRt:���+vȨ6�!H�9�#��CM�7���=��%��Ll�{#oYlN�b�ԑ�����\�
2�)ꕐ�4:z�lnUpyaq�i�_�i4�S�'�n�͈�G�.bh���X�^~��m�h�?�2�0޴�a�`M~�U��_�[%��e`@0�1��%�x�ڡo��0SңVN*�+����G��G�ǳW։��>��YU�5�]���N�Z�.gtߑ�NuI�0S�w����>螨�K���5x��6U��&|� k}&�+�R�`FuW��$*}W-2T�=��7��wo���a��J�^���i	BǄ@A���`��h@��@T,R��j���W�"�Ռ�����VD����bV/�@LnYp�ܽ�2�7����o$s@��ϋP%�ol���Ԗ���(��Q����_9>�I^v��@��2���Ϩ�	%�AR��F�# <D�!'"2;��GI���*&����,��4�@R2� 5����.,���Zz�"&eE��w� ���W0T�cPA�\$����>�9K$�N��]}(�����@s���ҏ�&l��������Kd�hD!L�]����G>�l�R��n��1QSw;H�[� b0�����sN{��V|i�=�����L\"��_��!'��Qz���U0���Bp��~�T:U��벟������#ԑІaʳ����27�UjNȸ�ͳ ��q�(��b��(��.�Gw�� �S�|��5����;^��$Si�Pr�-}�ʣ�]�7.{��/�<:��~��{:�f�Я-�M��̖�=��	��A�j�
��=�rZ�d�A{���
��b-M�m�?X�}������m*��B�L��%��D
�8F�g�����s�R�{_^����}Aݧ�`><Z���G�e����b��Ώ�0��ș�!gVƕw�-��v�W�a|�A�A�p	�BF���J�{���?I�c��/�'�y�d)�p��WӁ���8��;��y�Q�n�D�vNPc]�Dm����y_��Jj�+�0/)��)N������ wp-�u�N>��t?����>`؁�ecx�ʎ�������x ������T� ��?�f-��m���7��H�U�U��:� KixG�mv뇂Hr��}9�2�:C���=9X���3�s@���p��?��By�C�b;�����}�!�Eo��s��!��UCcr���N������Ss���*�
X���4�f�l��F]ѹU뛮}C�	�H�Ad�;��U�!�Mv��2%����2�\Lϵ%GJ�'�����0*��R	-z�$+��
�K�oG'a���}Z���Z)�V���l��m�']<1}��4]�y �(�vW�}���6�W-$�
-AE��^θ�H�������")�Z��&�|Ԭ�5�)�.��lH/L�P���o
<w���<�����ܝ<_о7�j���"��n�
���y�D��@Wׇt?��*��K�\�������0�[b��`n3Rr#�5��V����Lv	��������?,L���y�����+��3K+b{��!�f��㙓�6!��U�r�7�ZH"[��?�|0�ԋ��2�}΍H��*�l�!�� ��-��YXP��l#��ޖ38�'��N3y�Q�i�$��fh/ǐ�Al��#��wo�k�t��V_�<�T����~�)�]81��@
�D����1qqmTm0BmȩA��W�ԉ�h���}"��i&	�S3�=Dާ�ԝ�no��q��qd'�����!5l�A@�Uu����Oc'֕*㳷���{G�5�<�ʨ3f�P�-�S�}�����y�B^��)�*�
��m�N�g�&���� =���yw3�wR���5t=H����(Iͨ��O����;�N��Q�u�n]V���+��.{�~���t�aZc��Ņ�-2&IS��g䬍ߙ����Q��L�I�3�u`�ػ��ݭ:��XԊ�������HR�a8ԥ�xWs���U#�}$_���*-\)u�~!�h	���EE��0���<����n�i::�Rtht����߂c������!!��y����rq�	Oؾ�Z'~͵���nQt��|�����$������_9�!�~�l\��r�H�+������v� ��B��`�
vMB��b�%�h�"m;��'qu/B��va4�8�<�s�D�(�n��r��P8lES�{��e	��O)Z��h��9�y��Mn�gN!xUjI��r��=9�c�A:��d0�i����_1��4haJ��vvw��\GY���i�]�M�G�Wi̕4�]�P�a
����y�d���"�J�d�:HL�Bu@�r��= C�ktw��\��cAA�4a�o����L�����)�OZ���(����W��:`����t��������	z%����I=8�|�E�Ec
("\�n<�b�����yBV��ո�����G;p�A}d��E7�UI�֪o&[Y����DW!�{r��� ��),������e���ެ_�O���7���n���g��: ��5[PE�K��b�Mvo�\K����!ZY¨C��N�6�����B�����1%��"%ALF<3$Ӆ�ɖ�*7���%"�\b3����	��H��h�z�,(�L{�ͷ{K��P`>�=���ZƮd��w�i��I�fS�F�9�1)Yl�s޵�vz�&�93 ��$������Q_���z(�?R��qGTX�Y�C3�˸�]��D+�[t�v�"�2fUF�� ������r`f<��
~�=��O�����\�T����J�%�#j���IEˌ��o�Nn�!6ܝ�hk��J����xܛ�������m�Z@ґ�e�I�&������.|Sl5pa�;ۇ��+~e+����Q5'�T�EFb�q x=ͺ��c+�v�^}"�X�2�ۖ�k��C�K��?2�nH��%e@�(5�h�a���C�y��D�s����Bs�ss0ñk�~��O��˿� ��'��>x�r���H�"k�[� h���nU�o�	߫�b���`�f�*��ɵjŉ
1]���y�l���{�pK�.�ߟ��<��X[��']�c�NW��*���G�0T�<Ͳ���F�Ww��*�4���rV���ǭ�w,����	9�#u���-ƙ̀����������}����(��0�'*q3D���#�g��?='fhӖ�}]�B޺���C2�f�q$lk�eRy�r�������/=�^���e��?����S�+�[���Z�l|�ȌRn��D�{�Zt{~�P^�@�#Z��OŎ�Y��Qx0�ͣ~}:6)�~Y�|���<�'�����TxոOQ6R���T���[m���BA���[Ԑ-H́
J^��X<\��~$�c6��ɦR9d�:�
HZ��^r�*���<Y�	���-v���Pۛv�x��Ɋ�յj{)=�4>?�z�27�G)�k��MD���RuK�>T �$�Fb� ����@i�q؛7�p絤&R?c�4��&�5�����B:�{���,Pʸ�i���	&GC�ȂG��T�5�O�f,�<f �������Cƾ��]�G��Z�U�ˣ��~:�b�r���~d�d�K���7O�B�CB;�Y��w���yK�i�i�h%�	)x��yH���FIjr�d[P�o��;�H��q`��C�i߲��)��g��H�?C����㭌Qh�EO�X�ճ6��|�j��zڀ@�da��)��8�c#���t��6��,�I�4��N�ZJ�/��s�!�w���K�|�9��j��W8��m�r��& ���w[dQ(�j��#�Jj���WM��T�͔f��ש��Փ�ITjSqɕ���p�\ɂ+g�,��t-�2-h��[���h�Pt�6�i�E�H!�f�c~��nZո�Qq��t`��`o�Z��,Tɛ[�zم�ƣ@��w��N�u(�)��_�	�]���}�@�oL����	����`�6)]h����7ƢU�e,=r!��6��34lLr�tC�C����Z��)gK�����-1�H�����
�|�e�UL�a��s�&ɕjmO򪙛��Ն�K�g��E�x��ki�j������($��a�NS�o#�3�j��E�U�e��I���yj��8�׺R�Դ]/~m�	�s:L��H!%�(��?PB����81(�F2�1���P�LI-�<G�
�ކ�5r��Z�Z��s;}��v!k���9/8h!����]����vW�7��ڋ�X�A.�h�&J�Y��E���~�ڄ��g���O�p!��V�yI�i�*��1�]��]w?�� ��rq�̈Fh{�`Գ6-����X��I#�zr۔_d<���-�>�����h`p1,"�m)��Յ���s^}�(	u�]�L#��I=n���TG�9Q�����^ Oo�%.���@8��e��Ne�(�@r��d���)��T%����i�B���?��>qg�Kj79�IuBP��dU)*����'^X{�}�%=�1�<��F>�9���������"���3ؾΝ��}�{���LeO�r��ps�+2���K+����A�p�����L~3��w�&�^6py��y��R1���@� ���d���!(Z��%��C�[�TCJ`�hS�H�r�i&=�d��Ewf�|��Ӊk+�F��^�����U��
6ʤ7�Q;�̲S��xA�6�ȗ�r˪� F$�)��w��,;�oC�vln��uՃl�l.�+����m+/��3�~(����o,h?�t,�D 9�z�o���$(�BC��y?!�����Ƙ���)�1��@�P��a�A�?n���c�'�ݩ�l )���t��*#��K���&A�w�v�q�C�6wׅ��M{��k���^��J�Co���=��xl��)�Vj��:ި��kS�MdԈUdB:S��L_.�1 4RVk)ܕ���|s��Tin��喫�#ί�{Pw0��aa�|���..�X�`/�-�{��4m�/n�f��zG~c�K��E8H��\��ߛ!́��-F�<�e͕�y�_,T���#�5`��tZN7S�Q�'�7�D�����q��Ϝ�*�@��ri�-���;�,SgIT%�j0�ɺ�O�9���fsIvt}�����T�sJ�� ���}��=�i�B`MP��6+��1R��Ya�����N;��q�#�(�v�w��yΆ]�^��]m:���ﭲӻS%Xs�U��P�6Z�.h6��2H�#@�e�YP��aD|R}��(�W�Y�&P[����h�q�SGu�` �5q��_"b��-��F��%N�&��c7}�G�^��R�6*TX!�ۻgϫm�&�m#r�D#k9���|꫒1%I��o &����q'�IUN�zc�ٝӆ	
G�ԏ?$����n�Ng�IN�Vp��@XѶ�8����
�SI,�Ks�.������1���s���J��:�u?�p�_�)�F���۝v�?$�����G֒͛~�#����>!��&� ��n�Rh�Ji�/Ş�{��0��	���,U��Y?e1�1�<�V��<�����=��k�L[�6���,:���uK�̤U3&ykn���^�5j�'�D�~���vV�)�x���c���/��zS"��?)V��P\4�.�s"�w��<��sMIt}o�4%����2n��y2��nƙm�����|N��&`�B9��ҏ�]�Y�"�4I)������啔(1ٱ[[7�b��݇�Z���B�**�U�~>*����<�S�x	8��	'��*��K�k��f��fK �Y�>J5c��}{�ڽF��h"N�V�G�BC�qˋ���-WN�,O�*�;O��_�����3�v�7~�T4�VD�/�<��II�q������i\�����W���,"mm��#��hl7���b��xG�>7ܛ��;�Ѷ���ʑE|�sH��1\S��i)y]�;T��_7�@����L0+�����'0�y.N��
`&�\��ͅ}sLj���z�b��c� v�X���3ר>T�9	�&�ΛyM��^�E:�:�D|(�;	�3nI�*���C6�6¸
)Z�*.�F�%ݐ�2��sY�)M٢��ʶz�SĬ"Ic�DVSo�cF���~�}w��X�bQ:�:�/4\�B����a(m �5�f�r
A��,6��m�RH�Db�U�:�8m��#x-=�8�02���k�q89�^vb�k����CܕۙCO	�~h;o��N&�	�5NZA�0\�_:;�_�"6�3����qPHv�X*Π��o֓��� O����H��Ng�u��!�n��M=?Vu�U�����)(�5���#�Nv髢	"lz�^h�5��=����L�Vؔ�۩3����v<E��(*��myw�\��v��-RRAȖ�陘+T]��A��Ho�W�uA���可[�m��>�盷��f�q��,y^�cAA���֨�Υ��]�ޡ
ø�F�N��H\'u~T��7��F����T����&�Y�>��~�56e5<Lؘ�T�\ٓ!Co��qH8e>$�����q#�}�SJ%�[3ܔ�
Z�xXKm�@	��&OeO�&��4s3���2"^�l��XXF���`u�BR�[2;_o!(��t�C��=������`l��憫�^A2Ggx��#�����3��j&���:���'�B?�Pvrv2�!���Y�������x�� ���αÎ��j9���D��{�Nߥ& <ӱ��FM������V�J�)�O�eą��i�E��s�=w3�1 k"okR�(��Tҭ�tV:�@3���� �sbש�O,bj���k!6�U�M(�MF��l�S��'f������ul"�\��u=���v�.�.r3�~�bWe�-z�����]E��f-8kt�؄������w�]X�皋�*�sH]�+��U&ٳ�Z��財s�eŵD~�ζ��������ӰÆ���ߑ�\YL]'#=Shյ>����"!�4���2��;*�D5�Q����]m-�s�J׮B�=_jct&l��
�����oD�<��K�w�[|��g{m�J��[���=a���\�U[�>��&�V0���~=�f]3rv�6��5��/U�1�[;8c�D���f�����G&
�����Ƃ�;M����VFI0O%��>�H��-}H���ܘ�#��X�F����iߋ�A�	�Ͱ����C�͞k�x��ր�����Y����J�I��U��+��	9��Ai�zeV~���\�NwxVt��aB�*̒`�����%Z���Ȩ=������f���}ɓ�Wg*����+�;X0�b�㝢��7r%'늬��{#�u�:���g���<1`�U'j��i��<�@/��� �3k���@�/BhS~*)^�}2��$@�mS0���O#��SQ^!j=���یL����'Pj_�m�
���7�w&������S�$��e�*�ŭq�� Ĕ�n=��,��5
�%n��W.�؞���1q��,GgX+\����`��Q"j�Si�#mf�;ܮ+��*��s�Ü�.FR\�PL#��3 RU�:Cr�)R�F�A���(L��wU�<s��4�gft�!�'�����W��@����0�u�wgFٲ��:%lF�om�ht�"��1�Us�;�qґ�e�U�T >+��P�����Ó��>G�	�ٌ~1ү�$4��O��q=Đf�U�AajJ�T���ގ��ʓ�o�m��J�(o��m8�+ێx��1>"�2D[�%yL��=rxzt
`�\; ����Xl�q�zr(�'�Po���5ud -47dƤʌ�A|O��6wP5���)J��аϮy 0��B^�ڧ��e�U�͚B�?�@���o1�����FC˸+��VߜF���a�ͳ����9g�u7:+����Ga�W�.��߳��G�K�쉿R��c2��_��'mހ�;|��s迨�Ͼ�edɑ�V�����'���TЁ̜kQ�&S2�~N�
�/n�4h��}#S�����o�J_�XE*���ra��`�]���nN��9)ջs�������G��.@7��|y�z������ح�i�n����Y�c��Z�2ԙ��Oh8��hK��S��ls�R�q��nX������1���%�
��%ʦm�I4���d6E#���1ch�b]t����6�s:��*vC�|�~yM�
�=����|^�%3�n��kN��{��� ��<�n^[Wo�-��3�!�����2��V���s�|��V-_�L'v%��[9a�1�A��#��z��_��K��v;`2�K�Q�:�A,�q��H��o������9O�|yk�M)~Fj9%I��"&Z/�_���@� �ڣ	�'+l�0E��gѕ:����.JO%�����%3���N"���'����E�=���!��=,�sRxNp5���Km���2<�	�~I�p}*�k�&��Ǐz>7�S��n����"������.M�k(�l��\6� �~Q�Z�>�"�O��Մ�+W��V�QL�шv���
<���������q�<�M �_�)�4ȧŎƉ�|>��:RAV���!{յ�ơ"Y�F�N��~����K̿1tq�����`���A��J�H�ɥ��f�{mS��qb6��V]#�G
c.�n����&'KM;����ʵ�f�N�'��!�o�b�|艔��=U�w<����#�~�p���i"�M3�B���OQ�DB��*�;����L���r�q��11�G�xl��m���M�K�?`�xnFݫ�F����L�إJ��^:���)��1\��7��&���q[/�e��SMn�����ި؃W^'D�t��D����=7G�g7��mK5���Cw}���G|	i��'�x��N/̉��cR�������[IbY�({ z6v%�@����~䴌x5�~�o��S"6D�ɸ] ��I��b����4�8��w��gx�g��s,��F|!K��/Tp,/sD��5:��k�:�v�Ii9��9�OPZ��`��4y�Һ�<�a�@D8*q��&:fS��Y!�ͼ7�R0����{��k�$�X�m�4왰�v�08pB������Y�NZ�aV�����F��t��Uhb�.���d�D�[�6�M���l����D�.�FB�R'���p*hF�|����=D-<�����=5S�fJE�������^Ò�3�� ��eCC|o�^�`���),+h���<8���8H#:9�����X�'��f�l���"*��4����V���llwJ%���.�Z/
dY��id����0��LȀ$�t���K�ЀG�ć��A����z�YA�mɟ���驇.��Ï^�9�� ������Z�wQN�!�Q���ͬ�!���"��ר�X&���FmL�)}-�Px(�o���N��>�O@�q�?�+�P]�8���;_Qrm�p�D�K�.r�R2��a��5�Ȝ[�qR$,���!�5��h��~������&U)�Yo�����O����$Bk�+���
	�]G�2�A#���*hn�
������9w���\��G1g�<_9��(gZ�����dC��S�|�����v����v�h���mHd�sY�
!z��C���Wn-+W�s��Cϰ�^�P�ct��W$O�'@����LY�K:R=�(L��hDֆG��|�"_�E���aN!j�b��Uu�|S!v�D�^�����ǎx�ߩOVOH�^�<�b!�[s�2�����
��Э��֣���9�_�	�g�k����<�F��6�����6ե��j&�����.i�����dg۰0��#�^=��/�����%����-  J�����*���C�44i�2���]pF=2����2��Z����#+�w��]/�e}tNɻIơ�8���(��ʙ?d�W.�GT�;�3x��5<���XA�C����E4Xkn=2�WL�$~o2%�h����Y�f�I
��^w{�/�b�&���+�j��7@X���j6��;�"��9lA��H�@`dg���$��>�����,�4���w�Κ������YOin�AHl�:&/3�:ʀD���X<����V3r�I�gQdzt��ẓ	P���V�s�2���,����=��D�_�-��"0��Y;Cr!�5%D#
�[�y~�j}��y���9I$�� �OT���,/�wt<���<��mN�HU8^){�e
�}U<�nQ[�[�����7�=��A�'8&s�����|F�)�|�gS��3�q���7ؾ�f�g|�ڢH��'���r����7����(�,��UA�� s0��L��^���q`Y��9%�PHG_U����YSDUC\Ʌd�/�<��I=
�~Y��z���Ÿ���Hd���|D?��wc^-�݅&�M7���k�����j{���W�d�������|�c�}��=���8��2�}��G��I	�
�����`O��s� R��.��ݖlũ_�� �W���4j���1M,��H.fnc�5F����oQ�b�`bXhǳ�r]`k߱�䙅���$9_>�	5�_���V��ε�D��y�v�0'�P�����_��[
#������;44�O�X˴�X�yD��It�jS�څK��}�M�sՄ�^����'$�r��)��<tU4O����bZ$pݺ�M�;1d�S�N(d�,%�(��6Ѯ�?�nb�C�)���^��h�׳L!��"Q�CKq�l.�I�~�y�A����G���ׯB� nc��O��C�o	7_$:��}�x!}�gၱR�:��t���Gׄ�g�,�v����ЏL����(٬S�� m�{���x%)�_��v�m�X%����Si�rb�g��8�z�!KY�jh��bPZ��m��I]�}���ƌzľkP�?N�D��v��m(5�p��V5���j��e)X�3J��M�`d�7޽�m���(���GBJ~&�Umz�����ۅ����RW|�?6⡦E��N⼐���yY���%�(��/j��ޮ�#ok���4n&�8�.�r��R��|\@�#�����#��G��U"_�JX�}�vd���:��y���R9|H�v��a�h�:	�*!;�"|�Mv������Sm���Ta�c��r-�50��U�$Q+��N����D�f~�Ȏ=�0N_%V0 E�X��b��`�q�'��k���v.��%��3ݥ��;�4�����n�|e/
a���aN"�"P�r=�/�՞�����=↏(�8C@��_�+r�|x�{�U_$�H4T(t>���
�l)v�&��^p��8/]R��!2$�f����g�g�Y�(�����K�=�yp 5G:���s��7�x�����Dը�X�i�q*ЏF͉���'7O[H�[�����?o�Ǚ�{��"�V��Y�ts�J�B�R��_�6��@���,R���7���&X�8:V�K�O��5_
K�Rpr�I���$)�:�(2��?|1��y_T�f�6(�xf��y�����ڒs��Z�I!N)qX+�>��Oj�� �^��+d0Ң�u5#ʲz�J���v$�-�4s>~~]�4oՔ�W`
,*���:Gݮ}d D,y�,���b�7��&����"I�yp�7�)�Ce���kɞ��<��oo-/B�%H\x�m���!��=Q���N��;���5@w�ƄL�� Q����buE���.���6��۬���̩\���/�)�c<~�j����r
p;�Il�4�K���N������Y�}fe���76ۋ܆�Ց��Ȍ~#��]��C�ܽv�63�R�|�iE��D���j�#����FqV��6L���?x�G �%���fc>����g�{��G��EPeX�0�^F�+�
흑ۿ�zN�|���uY����`|��$\�@�4�����q��f��+��g��@�=}uِ�nb��d1��H�p��t㷮Ħo_�Ӑc'�dP̜� �+&xԹ�0�Q�DP�Jx��To�9D��2<��l�I�<0�3?]�8�G+�˩���r�ʭ�W�<{42�=�I�^M��V�����E�̎�M��+��6�q�//L�;eJ����������� �{>�x�ty���K_
������T�-#;`e�>�D��u{�2�".�_xzy��h��:��-c}9��i��U��i�X��<��v�4�(5� ���#9�2���>1�a����Xv�9��]�8�<'ӳ�k��Ft :����6#5�-DTv����茣��{ZL�҄�׺���{3���9ݸ�ɜM�-�6�@`N����r-E| L�_���d���N,�H"2y�����H3y��\�'k�{�a�+���Vy����s|G����T��$9��A���{2G�r����?��@R��͌kh�#�o��.%�l�C/�k�c!��uH��Rrģr6��6�R���s�x�iDX�Z΋�C�>Fk���aD�Y��u�Ű�=Jڋ{B`�8�c��S����M!;�E�f��H�֚;e�	�=+�@��ua�ǹ$��)u@m�bc0W-�Օ�F;u.%�s�9CQ�]΅u�����/��rv�^�UL��G2��k�@�D�JZ�	��tO�E~U>%�F�J<K���ѽ�vsce���7x͏2�ΧИmx5aO�h1%a(>A��D����:�F��ρ�Hxһ��F
]YՇ�\���e��������"^�Cm�,l��ԭRzu拦��#�j,��ѯNO�@:�<���;ǲSӋ�5½��?#�s�i��N��>j�oз̠~L��3�r�S��qBFp�W�˓�a�ޫmʙ �XtX�E�E������A��+#r�*�ʿ��y]�O�l�B�)����lB����ț�K�FR^'�����w1��S61H��vd>�~)�6�� �oSW�(Ê/k�\�x�Q�������m�� �K6�����ى�$�wxEKSg�0����N�DҜ~�q}��1���ގT�p�<C�$͗����<�b�4�=�K���C�ˆ��k�`���4 ,#p���򈔱`�֘H9�9�R���;�U�j��=Jm��{��s0bMꮇ��T��s�-,F��	���wE|��ۓW����h���Q�)�����
4��n0Ǯ�.���v�V���i9����D���jup&Z�ȑ9�dnk]��F�.��8�榤W��d�Gd�NR�k�m�L��Ů7
��"1H#ڶ"s6���KEj4J��)���yC+�$�_���i�J �6�`/��C&?�B����ާqe�.HCJWH�˨A�j�>�=V[�S��q[j��$:+yn�oF���\a��)��#�/ #g2.��9a�����F{����`���/�#��5��n��CG���X����#�h��0&˽�F�ٍ=g�&�Πs������D�
PN���x���X�&���.c����T/&|���F̪�C��֋l��lDC*��Z�%
�f�5�+����)��|f�]z�+�(���(�g��
Y~>�&ؑ*&PN��;c٨���٤��Z��];���)Q���^�V���@�i�Y�q�z�rCx+~z9ZѶ��@���7Y�S X�ߔ�a�9��]��I��3��Ӏ�n�%�|��|��`u:�׽���X��<`��Ѳ�i��W�	��J<�m5��JL�����Wda�}�����;��rx���(ʹW��޴4D~;�E/�b�LvU�e�[ا��GxО�l���Z�5�-[�=�޸���S�x`� �$�����M��z��&����D�6_��}�L�e�q�nV�	\#L�섦�$Txz,u�Ȏ�N��v��TM��`mb<@�TB��_��Ҝ�Y��p�����-���|�gs}�܀D�U{������Gqc�=� �R�M�;���"�`Q>�S�+@t��}�?�|��Va9D�B#�S���>ػ?5~��q:����7�Q��lr��	"*�.�z�4�;m=�:�����v��hqÖ��,+w�]S�JL��[;����n]��4(�Iz��Ng	F��x,v`[�͒N�q��Z֪��=��v�T�L/x���ѹr��Iv#I�4��ӼWI�Xb}��g�GV�?^��L('�u&�h�QF��U��"0��A8�s������R���M���	+4-�+�/���oB~T�&?~�	P�/Jp�eB
�����:PI�
�E_K/��{*s�㨘Ij�z��D�Wg�Œ�X�S��:�'��[}F��<�3�\�=���
�\�p���f���۳[QbR���$<lS��xBG}0b/#��u瘾��~Uᦧ���1�htR�������x&3��U�}�ZP��@b�Z2�t.�2k��@ֵ����笄����te��3��z��3����睈�1�~>��a�.�Y��i�7�
T��	�&/�/<h4;(o`��=�d�@i����v	�/�l�b�>Q�	xB�g���O�(k�#��H�����1�W��_x���6��J��w���r��ƍ@��q�t�-R���8,��C$�(�<��^��c�f�l�Gt���yߍ�I���e ��Pz�;4Y���5�mN�F�����nzO@�R=�~��:�Ds�����02?I�fa΂�,�md�(]l/����[�>w��L����#��1���%R/h��hn(Nv��5E��:�
bzt����!�m*����M��O{#�n���|��U\�H�z0������!�l��q�@�/f�B�|��$���|�V
 �p!�����&��/d�\B�W!9n��q5��T���;���䧦yn�gS
=�Lݵǭ+�!��J��JO�1�IL�w��󭖇��\'� �@5�̎��_�Z�ߨvxƽ���U�}%���28��k/��#Is�� gY����.���v|r�->��iw�mх�S�u,j�Srg-rʸ��zY�4N��x�n���>����~�<��u�J{1W���v{�N���.�����d���f~����eEGk�Hb�����?\x������G���(� �,͛�5���xk��W`���(����+�޽#�R�U���#x�X���\���MG�[iM�;1��d*�t��"ue�M���B��Q��ay� v�p��.�D���z	Z���� ��r�/�ɴ�tѫ�j`�ݯA�|N�5*����Q��+؀V|.�R�_�o�������뫣�]�L�*��O�������2+�@U-�=�c�]M�eE}0�E";�d^���uݪ!���1cR�7m�g�(E���}������"�r��Xp������!��ୠ��,}���-� �\]��'��3�X[0�"`�]�2kA�d6񮝘���Koej���pB�!$�Z-A%��FI�,9�%�!�k��S2m�3l$���3��*�	��H��k���"Ä6.��R�N F��k�1�$��5{��^����9W�>�����鿧3Cb�	���ޔ�KF�(5����V���Z�%��䡈��5�n!��z����t0����V�Ǎ�Pw��i�zmW���5z����ZW� ��D���FR�0�r���8�]ԟ�Zi���|�{��n3A�@�-.�m�)j�R��v[�v`�55��֐K����3����G/	H �\���z}Οވ,�wz�؎�o���pǃ�5�i� �q���z��!I�����*����S~�-��9��H0=C.�S
\�M@�.���z35�h�=��0��bw�8<�ÀV���2Й̘�λ���91�٣:4f�0��ޢ���dBK�\[��GsC����?���]�o' �>	CwXb�uTR� ����h´��$0�JZZ��C�%$����
u�D�E�N�ަ�@{%�
�^R��6�/�x
�|�$���e7��FJǅ&1b)8U\AU��mL�B(��w��7��+:g����f���ӡ�4������%tp�HT��y�.���	�x]g3u �{{��I-�c���^�W�LR�ؑ6��m�mj�	~�㢀AX�޿�e���D`y�/�� {5�vt
kv[/�kf(-�ID70P ��̘&�e懄Fz�#�dRN� �~2-o#hN����ep>f��Ov�9��&��ҌRE��+�dbL�c"V_��&��������x������.��)n��c+
��mM�n#I�=uֆ%�"�(2�y1H��j���[���:iϣ)�9BI�����p�c�&ճ\m�UI�
���ק�A	Ï'��i(���1�:GE�"z���׭�J� )�����<�V����4�跺&�[�G
�Q'�k�� �20���@O�l�?oo�~TA�5�Rq�On}i����8�D�����71d�v �b��2��h��A�h�
\�`�
�?}���-�{�}W� �T���d�~$��Mkm�K}�'��Zb1��TK�egI����Y�������x� ���.�R�Er0_G���粶a��^_�]����[��}Ap�z5(��B�A�q��������l��m�*��u��4#�����#3ؿ�O�	Kм������=���M�Ƶ�T$�-�SR[E"���V
iorNUAL1��'��校BR|V��L��?�խ ��ɌU��e1��Y�D2���N��ϓ��%®[﷠c�e4�𧀲��r����*?�t(g	�WaOYmy��|b$��2Fě���{�EN>O&�N�:`mg�ZO,c�D���s�N�iO7>{��٘V���W O1��Q����@�tD�<�ġ"[�y���a�%68ʮ&_�w����#b�U���W�c����ϫ,fҌ
����g�������0�����:�̂�� oM%8vk�@�̗�Y�V7�ޯ5�/h�[C�/Y�M+S�/����1w�8Y����!Idϝgc����oYP,C|Ie�ҽ���+�sh�$�@�п[�8�[�@�h�2x�3/��`��=P���:��� ]0���ړ�� ��YR|�c��� ��'v�aQ��Fi	���B",A�m����2L�sK7瀴A<����W�v:�VVc�wwf-l����Ro�
7�8z[�L<�.�?��u8�H���Hz~�	j<qV$´��M�ո��X�oy�"M4@�����������ú5|�I��"��359���j��]�D�#LP��
}���d#�gh�H��`�����t�{�O�uC����;gp�ࢮb��Vtے�l�I��~K�MeB��V���y*7���Q@rNuw�}�A -d���b �����ֶ��%�r�^_�T��t����P}IXwN<Gi��z^d��)�6f0P m)�q���G�&L�%M�,��2@��;��X��G�����T��|���
ԧ!6�:��{�pT�<�"Ӱ 
���ǋ�5��>]=�i�,��<w��s?��U"�>�b�#צC:������sg;Э�F��*������k3K��N��+�|��T'��Y�
�A*zj���S��җ\QTG�.�~��y���3�w����2K?o�ǂ��O��:S�]H����び}:9LQ���J	~U�:&�	� _�y�x�^Pvd?�ۿ���#7߱�)K�ǋ_�m��tw��u022.�B{`��J��U���e| ��BFҊRȆ�yr�����4�������H0�߾��'!?�2e-<R���k�WlԷ��zM��ǀ���� �����wFt�|ѡ/���a�E��������S��Z��t'��Xy�1�Ţd\dF��,�i��7v%@u��t�_��dKyV����*�FQ�!Z������q[�O��o����k:��i���~��1j�)��<7q��⊆��{	���n���]ca�ú-l��R�ND�i�aI��\n�h�fTX��ȞH�Ҏ�aA'u�|���C�I/`���)�Q�r�{W ;����|��[�gz�X�Lub�S_RQ.����{-�	�=��I�>��C������J��	������u��n�5c��9�Gu�� ��/�1��LqH��3�KQ�Oz樕��'��ʏ;�?��n�̰m|�]։�u�U�3G\M٩�Vt�])���U���U�:Omzp��Pg	��[�v\���o�m7��n��Jn	.��xfj~�z9 dh��G�`��Bԃ�>���O�f��3�0f)*������ҩn$��
��	�sQy�γB���*�&�=���-Ā4>�h�#��B�����vp����_�K��4M�Y�<�LO�KfB>�:h� ޸"]Iσ40|X�p�#汀����j�*�\�1S�����z)�E��G�3*�g�s�
���p/�V�THG�����r�H����+�A�<����%	6��
�ZO��@��|}�ҥ����_<<W�5�{x��T
����e0_	{ ΉDkw�@�-�6�7���Ֆ8U��\ٸP���'�kf�P_�t����#u���	o�0��Msu��+������~X�5�ڇy��I2���aA��l��[}U��B�|Ǵ4�&��s�~$�sN�@��f���o���V<Cz�B�۶??x���X#�,H@]�hؚo��Ч6��'ϻ:�<�65�'�1����W5��x{leMZ j��NpR�I�K�a�L7�2���
v�/t���iF���k����#�$)��H�^�7��F	��ќ�X��6�����:��ӗ��wj<��
G��}��D�޺k@ŉ�n&i��2<��9�^vY�W�,�'��2�}�+�h2�\�y�p�&3|�5?�i��yX'��=9���h�c	�n�!���?ؐo���j^��Y;�e1�l�j�zA�8[��6�����$P��h��X�/��|�	-����Z�&��Ћ �0�����EՀ�I1-ӄ�  A��Aud�� �d^`�%ڟp=I��v�4��+W;��|N޸�w��l��w����,�J�~̇ϐ�z�:A�N�p��_����Y]�"eO%ة�F�#S��LJ̦ԖnLWb��iؕA�er�oWG.�1�
���g٩B�m�E��y��FmL)�@̡lGxc��5��5gU_>�MJ�u�G���߯֞�����0�BpoC_��s"�A;��TO��:#e��?���gҚgD�3_��ق6f
�쀛=x�Yخ��p��/�l@�)��m(T��b�z��u
Q�!��l_��۲�
#k#6d�*]w�}� �񋳪��추A8_/����A�	a�T�6�Z�O@?#�Q�_$G��Lmў�;�9�ɗҥ�e�Od��М������c>�`go(g������������c�ha�JA�~	��;�Z{!L�4��^�����Nk^��9����٤Ϝ��q	�p��0
��8������4�i����S��X�ε��#Y!W��e��=Rƾ�c3�VKVc�E�����UG	Q�2�j�"��+@cn7��p�VfŊ��f���F�p��H��
2�<	�Q��qث����w*J���XK �O��2�v7�m��z�崛�dBM���f�R�UHOWR8a�K6r��ҍ�������[[ =�.Q�rPTJگ�i�0b�7��MlP�)��^��7���~?��������e��sM;�w�N��L{ՑV���K_P&��^-L�Ԛ���J��sԂY��U�&�͘(�.h`8?6��G��j��9R�c�����ǫ�_���k�nϐ|���Eؠ׎���a����"�w�w��a�@�X���.�)�����JL�����V�=��D��UK�t)��V[�.�+�6r�p�b&��