��/  ���#[��}/۷H.?y�H����Rx���R�}�����V�!f�n7'� Y�%���i��uxc���.�∶���=�{jE�=�$a�����U������_f�_@C[���B�}3Upj�d��c�K4��u�̿K�WM����P��n���a�ƕ��.�2_"�jGT�˚J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&ܝX,`c������ߔ�ꏹö�h��&=bQ8�[lYXDA�f�`n���O� ը�fN��@A�M�5�l�m���P")�j�=�"d��e�����%�}F��$�xVFhk*M�Y��0B��5��>��Eॄ�����+��t��Bh���Ld�u'*�j*���xn��t��`���ˌ�*��}�fT���Ց���D}�RI��Cu�����(� I
���kt��!E�� 4��fN_g!�����݆vo�J����
��sP�ݕ=�z�E�5pc�{�w�f���[�|W 6���.���l�&�ii4�񰠛��� }Pk�g�,aCj) �9�L;��&ͼFʢ���e�0JjEB�C��L��I���6�D���j�.)E�ʂ^.��Kp�,E�7JTt�����c5����#_�VW��������"������bUu��:����uPK�]4���Cp������P܎o�X�Dr�bF	�b��D��0�DJh�}�f��x�}��L���M��-�%U��G���L�hDx�^�kp�1�&�4�� �C�����&"����o�Z�p�v4����A�8q �����E���� XjG����s���N��+~t>J����s����Ͼł�|}d�g�S&�s��y�l�btʃ�����f)��ہ�F��)�K
ᩢ@\�����|z��y!���̞B��`��A��"�<����ie'��� �.�#f#(����>�1�M�f�R����abU�D:�ɧU;�W}؟A�X�8�̅����?F� �#t*\MaS�4L�-�����oF�},t�H�D��&�����g�4���Y]R@�wB� YԚ�������.�3���!q�<ᵴ͜Atg�ӿ�ZX���r�Q[��K^��Q^�tL��3G\g��|Pb}�׎ɮ��4�6�Z HX0�!e��/���)}�i�r+�6�p':�6V��\�Q����^0U�Wtw_3�J�#雔5�e��o|%u�[O�x�4Ʊ���=�x�@V��G2)#�;;��FF�	�p���x����kb���
N�r��xpM��(��b����X,�U��c|�Mȫj-�%���|���+>;q�{/�QaG���/f�{�b� �6��**���tIf݌�?\� �)�,-K��z�D�)X��H'��CiRtmY:p�n.�K��
`�VːH*��L�B �����>��r�JRӺ�{ ��\/MҪ T�/�Y����i&�����S�R�3��Wp[�@�10��T|Kղ��r� ʈ�v�s���^���!^h�`N����f�h0~\,��YWpѿ�%^3Hh�+λ��-)6�0辽e�I��ɍ`L7�d�?�X�=|�!���	�o=r��v�LK�EBM��zF�N�Ds_|-EC9������K�`/4ME���D�|R��C���T�"��U��gF�.�#���X{�� H�a�ucV�&�$J[��sQ���#s�9����].�~���0�*��+#lr�B̽`��)�' Q�U0$�Xei[�a��5drY�^y�{�>�G�=��C���9N����[��'��J�a���#I~DI�O��<���߳�����hz-�Pg������,�μ����;`�a~�*�є�`2�B��A�ǰ��Fψg��Z�{و	!�UR|�'��{��-�w�X����.v{�cH��W%��eaC�H����2��'Q���"�j�+�Ӗ��Z�	�UQ���{K���
%���Ɛ�z�D5h�Y��9֗N��,�@�'�����u�{�N.��e�ӲY�^R�5/�����{���OK��>8(W��y�	v�~+̂!���m��1Y���ǂ��rdp�'d�_��g0��Y{�e��1)W�r�E�D]S�Y0�(v"��'܎k9<*Q_���;��w�8 ��-S�-�B�3��O��%�JWߪMl����ͤ��r��5Q�kX���R1�Q�U�b^�x���j&���X0�`J��@l�[�E����v�p�b��d6v�0)aӃ#��={b����{�0h?X;��B�%C�SxwfϤ��C�۟X��`��و���З��i����51��
�D	�MŸAƴ��6�%�:@���A�S��&�;��M:'�<��e�/�<�\5��-,Q�$���8�������A�}�H�4�?at�l���x�j�>{W3����$�ນ�����W���˝
�\��,P�p��O� � 8��Y}
��5$���3����rW�Bh�t�mk�=[56w��eW�`�Bs/ӑ�sբ��c!a��j�v��d�~R�[�5M� �V�AUϳ��,�Fe Ɋw�D�Kk1f��	�{����2ԷG]a~Ҍ���ߢ�φ����Q�`�AtKJ��8���31�&�����6\���\�Y��tDd~��!���3R������_��N�U|�An�e۝�|�؆�}��-��e�0�3�$� se�a��a��ڛ��|C/�H_���_Bk���L��$�	.�f�}f�2���D���,��Z��#��J����^AotO��u9�v�E� ����*W~�Km޳iW���g�TfS��+n!���)�h{f����wE`��cQv�$�V����H���]��޴i+�ۖc�[�w=��>c�q�E�W0M�B��D��!���{�����=�r(�/VwHFx:Z��vL2��s�T���TW���1E�5}3W����V�A	m
��B�����,K/
��KTZ��˱%�|~�I*HȘ��Qı~��e�; tʘj��SU�V����i&E!�Tg�W��Լf�y��0�U��	$�� �1�HMޒ!μ�5S_���F�y�bT��aFɃ�����s^����VCve#�P��SD �4��|зvXQw���AEKAԵ�p1V����-��ďH����E�����"<�G��m4iz�'](	 �"["Lܡu(�j�a�EE��<�,�#|t���Ej��^w���*v(��<�C���{r�B)5�;Ǘ%K`��cTh��⁝�󊽦�ʺ��'Be*�o�Sj�|u/fZ���/�
 <(<}^��s�F �_�B���/�n�U58kw;vl��^�Ɇ6�\���p�d����E2>����)d����Q��gO�E�]��
j��%h�oG��ܸ�ic��u�#]���Ϩ|�wwsS%ނ+���:
9��ł����Z��e*�>��vsbF��������ae͋l/���7jW����{�²9�3��(�t$dsf�%�T7(��{���};]8��0��v���Kv�(�s-=(�����]�]�<��S��UZ6~~��o=1 璼�=��o"��w%Z��!侂;�^�q��{ �l{#�Wgx��~��(\��ښ������cn��O`0�`e;��%X�5	P?�Ta���2��sl�b�����ᜐ{�S�+����`�'���N%&��W��;��Kن��T�Q:��C?�VJ}�^����T�M��r���)�楱��53����Ԥ/��ijn^U�Kw�S1��u���2{C�3�m}g�+��tW�_��� �]���;�%W8���b�l_�`�	i��(_�p��MN��S 㠝�-`:��&\�ʔWf��E.h���f/\��Q�D� t���pFlf�z��U.㹃�-Sc�Oq�bR�P��I����j�����3,FHH���i#]�E93���|BH�l�zY����ޤ^�(t5�B/�\o�qs�#ɒB'jw��d�"i<�,�$+���]��[jr�t�M, ,�3���͂v�9�R�$�>iñoD����r��n�p����<(�%��[����B��@E�wq�M@&�~{�"�+��.N�� ����h�3�Ⱦ�@L��&ש����_{}�7�;3�JY4���UVV��B	�[1����9}�I9Yx�Kl+Bqܔl9N&�(c��Z\�t� V�=�?�N]�s4�,[�!J�=��{��϶'��g��G�9�������� u3>��~7���ۙ�v�:��F��b�d�q ;�.���[鵺�D��%�<�+����.�l�-O>4�x-�������Y��K�-�{hs�T��Ӟ��c���8���:��ֻ������m:#J��UV.~ɫp�����km����P�k	� ��ϾgZB��,���?�[G�\��<˘=���a��Q�qBт�dc�3�Ь65�L��䎙7*�X�5;g˫���D���Z��"�A���Ȳ)8�e*�[�, �K���#���^f���i���"���6�ܩE�32��ɷ����_�B��Zˌ�}$W���^���Ɩ�q���OuY���B�Y����`YQBD_���K�)�"�rb:��+�Q'v����.��hNc��}�� �䀪
�͑_@G�ۦ�AD��&��'�5�U�V��b��xF߇F�aӄ8Dw,�B�0}�iז
��\Y����0�oaE3)z��`��w���^��R�]$4�~^(u+-������*	��>\W$�1L�-=�t�#ɞ�+2%�l��Ȏ��{�����)�)V6�Z�Yѻ�R�V)��H��^�}�� kS�h�����Y�k�C����A�O#mq!P��>geK��uC��Z[N}S 6:V��@.���*�A�x{|uZ�77w:UM���q\�e�{��3ŕF4ۖP��Ew��V�i!�I��E���$�Í��ꍯŇ~le���_h�b ����� ���ߺs�K�u��XWIN�ۨ�k@�����k{ux?O��+�rK�w�ئ�ٖk\��S�xMH���X�D���/�YѰN�$	h�U�Y��6:��rE_�'՟۞1�6&�
 �i��K��� �gtS����lb���ѩ��lD�]w�����3yUb�z4�7�y�@g�h�u/K�GX&�2Հ�٘��HK�>*��j��lۑ���̜{����2�좨Kk�����s��{vl(Ʋ���+��?�-�	��d5��M����I�aO��v".ߨ������)�^�EI��=Pcy�޻�_�D?��b����Ŀ�S������J�U�\���7Vt���
\M�Z�,b)O�]+����`�g�r�h�b�P8}8;��-˲0Y�8��޵�p0��p83*qO�Ț�,O�n�m����I{�'����"IR���&0�#����I���X��%/fOӵ����w߫��&��rK�T.r�a��d�,xzg���*{�s�yx2<�dzjP'�S�T�~��|YG��BO��kYd��7��r��z�*��ȣ��1��'Ѷ��l.���mfw��H�s
 jQڽ�9��)��6�{�s���b>�рc��G�n���Zi7�sB��+��{�㞿z�h�T�5X�!������#��E4-�Cz�B&;5\��j�ߡ��8���P���g4��f���v�w�?h��AKB�^x$�����)�i9�ȴS��$ÁY��1S��zRg�06,����7������'�c��/�t�S�8��9>ۼ��nV�E�} ��W!��m?_J(�(����v�gLΐ,��B����?�Ze�J���w}����+�����wm�&Zv�{zMt���f�T�'�CƐ�@���ٳ}13���z���}'���h�[zs7�E4 ���n~�a�d����m���!ق�P��!D����Pw��ْ�z]p],h�E��(���K}�L� �kO���N��}q�(U;����	�~n���)�ʞCd!����m/�)�z�OV"�Ө��~�;c�V�'u�͵E��W",Mٔ�-�����De�@p����#|@��w]R�t͓��pbb�J�n(T	�����
\aZ�?`R�l�xl���"9 κ���J�h�Qg�@d�Ƙ�7��p�����_�+Ki^��q�[z���z_1n_�}7�~hZ1i<p
���&�q�0֦�����'�7�hsXv�:y���5RJw_�Gx�TgI��.�ؿ��uGeA�!AL��[���I��>���['G�����N ���w�U��W�y�:�u���Į6]�ق�'��#X>�^�;��;M�O}X�^��i���&8Vb���Zq�XY.;�5�?�-�++hϵz��5�����Ƒ�Ut�T=�p��ȇ����Ş��6��X���$��&��p5��K�&�+1&�y�;�=&��b�=���?�D�A�$̤�f\]��J2<Yb�j��Hb��!�[����^&�`eOU��|Qum��7Dl����uEr�E��m�0^�;]D�i�>C�jk��� �� ��mmb=M����S9����4�kDz��m��m��%M(U?>!��FK���I�¾Y�;���t�\P�*n��?�s���3&`�av��o�v����o3.Y:�)?�w��;F�����c(KMM��+@C��$�N2�i���_�S�j'E������,LX�=�4�����Ţ#��Ƅ�{^�"W��Z�<�8�l)�bv�ޯ�BL�NL���e9_J3������k�Ҫo�\���E}\�#[.��l�0]b���%Pғo0�����Z�������[۝&Qk�-19�N�*��нӹ��VQ5~Z�c�sb���+y՛=�T��A{�ך]�~r<�_+��
T;��Y)/������'�U�3���7x�_��r{(#�����?��޸�b?낺g7�ӿq���P������<�JOx��wp�ÉɄb�k!6�����z%'�:*�\v���Z��� �5�:|�8��aHA��ؓw��s]�5g`�_ds��j%1���P��,j�}�l`kZ�-H�l���ا!�ަ��kU/�BY�%㌔�q�'-���*��scD���A���=ޣ4D����A��S���f%���#h8�����xBW�>ۇ1v�����H��3�Z����:2��	��RKG�"�6�f��e�#�D�gٛUnvs���ͦ��BMV��n���cG�Ckfڹ� �T���TP��_����'k�{~��ɸd��ro���CUa�j^�N/D�
��(P����+��\�0��ՉD�cn	f��0\Å�Ē�|�B����"��Ǝ������W~>4!�62tNR~F^.�t+��^����x0��Q�AZO�:��9+�UlY��-un�����$`,�N������m��ի�%7rҲ�*ѵ���Ka������J���X�L�;. �2�~��0^��}<v*���v��x�Y=·Гܕ��������?�z7��ߚ�6f���&	P��w9	N�ֵ��]���D��LἩ 0�5!LfF\�����͞W�GR4�n�a��<�Iת%��>v:/��Y�F�}ql���PK�'Zg�ag�7W1����>���t�B*閍��7�w����(D�,M]vv�벱S����K��\K��o��š���	��Ҵr���s�h��`�랣��w����'��Ny`� d'�1�2��:X��oӘ!��,D�vm�Ǥ�vˆ��A����T	Rg8[��2��ؽ��@�^T`{���)t��Ae��)����\�Q/��?�0NS�d3��"�qv<b�J�0�!,�>�p����Ti`fL��4-w%i*",&/.�~��x�W�>�_�4(ϴ �J)��������.�G�tƁ�t��+�["d{�mR�-��C=��5#�s��� ?��pՊ�k�M�/At�㜺����bNQƴ��!%Yb�尶q��Tbd�u#Q�7;N߆r[��I�G������[�?ܥ�莹�|�����d�t
�[�܋-�1�� �-S.̑6��x��-en�	��?WQ�$���*ywW�-���>�	�cW;)�Ud{��G�Ѩ�)/�#�{�� HrX�̃�W�e�Qtm�3A,�V�z�K:S7-8R����j�ht��|��;[�����c�1]�
��g%tr���6y�8�U��Uׁnp���*���W��Z'��Je��'[�g}�ԙ֢K/G%_5��=�([zl�M��C�F�L��%�ssk' �\���>6��!X��f��B��vU����z���u]�y��(���VBڣ��B�|�<�S�?\�b7����v)�gJ`�JQ0I� �P�&�͙z�ƺ0I��8�琦��:#�\��ZI�zD-V���8#�x334Un�3���a�7�ͮxx)ߠyK��)�v.�<����O����i��	Sʚ�����og*Ź5-��K%��l�g�����]��(���{� tU�k�C�"wY� P�j�-e���P݇���#*�6�qo��٣H����ϡ:��P�
P��w�7�@���n�a�Ao]���s+�(MN��$s�������G?��Yun.8��ܺ'Wђ��\���$Z_j7�v M��e��f|��-|.d'�F7ڲ���=I��$���|�����W���h+��ʘ����� ([=E����؇�Ew���X�m���{����h��L���/���P[�,N ��ˡ{�V�����QY�gld���F�[�� .��j50�s�`��7,@R�7=�(�k�d�rt��cD#�7�=#2xK�
ئ�$�2��"��~
2kӶgM�;qJ���hy�q�^����#����p��Ƣ��Bn�\�cr���gjbp��[�&�B��w�BxJ�쨏��|�GHm�><���@������������Gd�%쳀�7�����왘�/Ov$ug�?Q���q/X**�3Тw��`^���v��̗m ��7�	�d��\����է;˨N��^K�	 ����li�-w�:��o��=a^�W?���$�,�_���=��%�p�Р
�rS������˦HG��"��0zex������?ɑm�paVH~ZUE�yUTG&����� r�i�Ay0iK��)�[Kz2{>��6ڋ�d�=�t����W'TWS�2�����{���;���t Fʭ����-7l^;���
�̚�Ѷ����c= �5R����S\s�5���(՛�W<��s��*�m�'<9�|��=v�ϗٗSV�s�R�]{��u1��^)�>z�:q� hC������~�f���cO!��I�9�
ϯ��;�ybq�t�]�n��m��P:��kW��}.���ZgԲ�2���<���,�;�=t�q���Sf�.ME��?]�u������L��e�3�bd�w�=�ga_��!��"un�B�&$�z�z4���a���$�k��׹�t?ٜ��%�6B�Rv���a���fk� ��Y���d��x�af]�:�n�K�Gs�z�O���d�3�^B�zl���7\@`̟$����GBfG�٫�y��;M�l�㟱�湨�6�s(/1�]��f�xE�\�r�i��?r2�и)1��\G��n��dt-�5>o8rq1�>s#���=�j	�w������K��C�%g�s�jN]�{���i8�TZ�F��P���!ї�2U�0�0e������J�����Ig֧����t:5��=����kD��_��ꐴ�N��F�:�%���u׋����X~������E�s�̰�g�ߕ�RH�
J%�ⴢ�6���i����wDrЙ�ĕ��=��Kҍ*������w9�"��VamW�uѶC�ߓtܕ�������n_:�u�c|s�h|ls�0Ho�/	f�H��iۗ>�7�ɿvq�4��߯��W��V"ޙ����K���4}��Sl�A����Ga�Oc���1t�{u^G��$Œ~�x�.7���Q ƐVU��D��%|�v�8L�PK���gW~*a})�GU8���Z+�4�X�L�M ����l>����?��J+k� +�f�EFh�z�ܯJ��@Q]����t�vx~�pF�+R2I�hu�}R�
�_ε9&�0�8���,�4@t�It���ř��u�J���wGЏ��0��a��"d@��P�B�:���ǫ" �f�����sV��u�&�Z�U�����߿U��Ð��CH涷C,k}�b�bE���~L���O��=�h�GX98e2�nJ^<�}��H9��=<H}�$�%��"8���?]6�1E�J�I��x�]M;�TP���YʐV�/ ,��J�m>+w޽(��*�(������ұgM6(�z��<6���׭d�X�yK�^��g�"�|��exX�l6veӐ/���^�L(8���!�Y��@Et?B$�����j+�d(���ؽAyVH}/SΈ�@��}�s/�4*>���En�8�挵��4�F`�{E~�<��M��6�E�*vz	.C|#<a+���SBm��_47Φ��}[��$".��-��@�I ���W�bO�?���I��bX����=�;�I{ v�w6�"�%+~UT��JƢ]n�Ʊ��"���p�K~�;�=_��}R�=���4��$.��-�߉&F���M]��HO=�� w������e7��38�`(�c��ZHx�oT�����`5vW����`%�-~ǫ�x����'P��2Zx�h�O��c�lt��U�y��3���	�Q�B���Q;��(!GH&g�i-���Y�}t��,)Q�52���J�e.�{JZ9o&%�Ĩ�[H����B?��KA$ U@��
P8���E���R��j�����?/)t#�2���LtY��F�� u��i�hM�]P�ܥ���P�_��֦�\�	���-�5���˧r?Nӝ+`���ǎ}�"/���p"k�,��'�|����������.�1B˾asB>�c1�1�T��~/Xn_�LT��5I��>�F��ν�XG�z#�R��.r�-q�s�<�25=G�/��%4)�H���*�h����C�>�sY	�?�%��ޮ�*ۋ���c1�w�Ȯ9��Lv1�/���r�F0�0��FBn�{�z��4�jȟ��0߱�A�V�\��rB��`_ǜF}c�$��t���|�oZ�9j;_�	-�@L
��s�[�:�C�MJls����1w�ӗ��f�A.���80�x ���2q���>�y�R��84@�V"�yo<奂�R�y�"f��E�Lƾ�0zpy�Qt����;|���}-��Ax�yQ��.q˙�e����,�zI0H�&�BR�kpN�Aҭ�o/iDЏ��I�^�R$����:�����!p����{���k�J+�A	BgE�����^^cm�����b�e��� !�oJ�`��/��؛@}�&��uGi�/V"�ck#����OA�r�Wvm�����g�D ���3jς���K ���
I�3�����  ����cz������br^R�mr��7��s)�sf��c�es��<�rJvt>:�X�.�q��h$@@��ݭ�Y����.��$�,��g��b�'�vR	�}+���U��Iw���A֔=��-�PHdZ�r�I��.~T\���Rז�	��f�D��(�����U<�̢�β������l,����i�����ЁYih\�3��@}&ް{�o5�kOsʍ�0��w2�@̯����úO�-;$c�m�V�u�5��6��c6��	�;p^��� ��c�QF�V�P*��Y:�n������c4��b��<��?���>�TMD� ]�GD��N�ٌb*1k��oۤ�Y��u"j�/a�9�;���4�R�g��ׁi�2dI��m(Jv�������s?pA~�1���1�lPG�4v�003tO�f��7�>}�ĩ*^3��oa��E�ft��o�"�! �t���e��b����5�V��\�!��`G {��t�\��h�"���S�cܭ�e>_�8����@��EV��n ҏpCPcZ�\C�� �S^�U?g��|Q�:�k��}?�m��4�H�'������?f�<qG��Q��7�c�m�]��9SHmFr���&x5�i�>W����cy�\8�H����fl��RtS�U��T�~"#E���!�J��:i�nJ�� Ns�!�
���b=��qt{G�9��տހF*}��V=��^���(�A�0����l�~Ԫ*͍&�-n+�/��	.��Y3�q"0�f�{�6��z��R[�e��Ef�G[~�J>��le��P�����Γ�8]5�!�7(��ϝ`.��I0clW�	�5�|6۽9�cWz.n�(X76���GVsNt��t��E(���,�iڪ�D~�� ��g���������=E��$4	;F$�e����u�,p�&�ށ�J31F��˖�ˑ3$Xe�@ڒm})�O㬛��
�� ��<�������?��B,,���j�"2SΈu7K�u�.��&�]Zx#ZG�+��_�������@ڦ��kV��g��4������;�!u4���C3��z�m������H�4+��N�\T����:$_+�0�&3�6������c�bs�!@���y������ '\�Y��k޵)��,�O8�h�Ϭp�DڹuY�I�&��2�0�u��q�&m�2��`���t���P48�_�Ni��k����Ưw%gK-�.�Z�c�(�z��F�K�T!���O���p��;z�0�F����q��nM#rvR�=�E~��z_�&��`�:�AQ��DP1�f��]�[��mu�I1���ڠ��`�(&|��"Qy��B�I��x���E��������(�.,���F���L!%^�mæ�������u )�3�t�/��F��v*�,���x����k�Zx׳s{�|���1�卋8'��'Y�}�����j�]L��E�v�:*���ŝm ���׵�ۗ\<s�Yh�L�'�"-���ޔ@�n ���Aؑ�΃�|�M(H�u&����)d͟�;����kl�%#�p��_<��TH(l���|ٞ^+�K�D^�f�
YJ�[��%+p=w_���P�1������R�Q�y���H�|^�'p�|2ε�\#�MAs���m/@�U:��������n�\.hv!�cR�������f�kT���/��9�#�{��u���ˉs#%N>:\�q�G֯����3-�`�$<:�r4h�*4��&�_�	��04��VF�õ��`�}�wC���d�66���ˠ}�$6�p�'�k��"c�6;��z�S���b~aW��QY�������Y�8���X<����$6 aV@m�����@i窢�`���;�*kX�Zm�`�*2w�Є^��R���������F%+P.�.s1�+�8~p�1i�9c��gT�F[���J�d�F��������g3'�"�,Π��_.~�>H�l_[%�Dz����ce͔��H�S�S[�4+DhV���J2!Y������ ��;0V������@�x�Z.�կ�;+'YM�ߙ��Λ�������|׃�-	B��G� Dª�~�T�ѭ����[ׅ�~��z3s^�\�[K}9Y�J'�ܡ:Gہ��&���ƨ���sD�"F$���?J�.��t�|Mҕ�/>3ߚ���'�i��b��b�&J�*��c�n{�_EPj�$O�(�4��'�`'���(��5�\??�y�]pJΥ��X�Y�Tl��&L�'UDl�໌���<�Lq��op�@��zC.�̅oq����D���fP��|y�8��JZ��ߚe!M�m�<r�ت�XQ+9Y肂!���^O5�=���0P����j�5<�S��m��l�3~jd�,2��C;��$�q�)�e(Uc�$�����?w9��(��[6��A�O��eo�H���)\���1�+�z],*��^v����gz'L�8�.�b'���M���Y_��1}��؝�|#;��:?��"T�{x 7�E�r����ժ����4�G�ىm��s�`������8�����_R���4p:7��e�� 'BA~<)�+P'�����"�9pe��d�������-�#������U���z�k��~⥧ztz��]��j��4�%�Z�z���9Ms�#�)԰�A�����3���W��`OM����HKvN��d��S��X9�lq��U�3�m���k�IL�����|�N#q'G[nX��� ��U�e��8��Q����&V�LFS���ڼU���ǝJ ��Нi��_���1>>8���NF(X
$��A"�C&4��L�%��;�E�9�/tg�r-�S������W;�[:��g��{ nr���b�%��\B+��Q����|d*	N)i��$	W�_��`�
����eĴ���F���9B����D�	�RYyjSQ��43�pdҧZ�~����Lv�u	�w��	���
�'"USs;U�f���Z���z�r���X�%�2��1Ohn������8�(��!&,Is�0�j�]�A���eV�%O����v�����I����ݤ�B�Dl(�����F�� Y��8SX�!�Z4*ч%3�f_���z:��-�{is�.Hw`B��i�C��:��^ uّ����4�2me6�]�t4n�_wc
�^����� >����5+���S[����a�4�$UH`ǿq�?��{z�B��Z��Vv����¦,Sg�U�C゘=�۰K�r ⲷ4�}��|���:�������QHw�D���m�4o�y[]3�#�X-1���q��ѩ{�	A�ocQV�q�d��_� �y��ʥ]0� �Ȋg�!Ĝ�gV�w��|��1�(��; � �_'�7��_Қ�S��?�.D��+2@R����R��e��F�O2Z��F��t��Xa銻�5��&��{�����1���1��Q��"�T6GO�\�$9�l�l����;��^��ͦ��B�{��9G� '�FU�gw*E��fcd���9K����8�A5"M/�%0�Z��R��ų�:5�RVJk��oh˵A��HJ�=�9��B����KsN8��jo���)_q���_d<?�ƿ��<�*T54��+�T�C�ީg�z@Ũi.������ �!�C���#7C� h�*s��v ����iv^/�U�bKY�%(�� 
�1R��,�*L����ˍ��پP��T�O1�w�d�^cA�cU�ӣ]NK���d�!8��� áF(��i�����-'hX?�~O?��w�ΰM�@g� �	�"��.�S0 |�Lcx�V��s9�:� ���ͧe�p`L��S�����Ź�vB�m.�c4�[,a�gY��������&ܬlr�P�w�9���M��p_��D���\z���_��>�,Vi���r*��2o�BY<{r긌�����r�A�m�&ߖ�L;N(�J�)�7<����bRZy��K"�*�i�=�9;ZT|]d L\���)�ׯ"����HE��>���[�v�����ZC����f4 ����b��� z&��(_�t����S� u.��d-]Q׍�OJ+3��U��}�
�4������4�}($;s��`=��*�Kͼ��b�&�&��.�{�
ϙ{���HI�X�O��P��ƣv��u\e�ȸH�E[<-Q=�*�ַ��zz�����$ĥ���!i.mLf�ۄ��
I/_5�왷W���l�	^V��O��Fvl�',K��͢Q�{�/��B:����`�4��5:�LpD%��:��� � b=u�J	ہ ��[k`��e����XT��O]��ݸ�`E������IH��+]�}��v��7Ӻ�P93^��@���������:��qr�@�?,g�O�/E*���j���tT+<�8�`r�p�PM�2�uR��u/�����NZ��S��6@��*�u(���u�
$�~��2C�V���[�f%�VD�����9)՚d4|����PT�O!K'�y,:�t��a����G��t�}2]�ۈ�0���C�	,��Jq8�� A�?Y#��U��8�;O�`��S���x�N��ƽ�C-u����J������.���0�p��>�WBNW�Ѭ<�g��/.=�P�r8����j��M��Q�*��ZC�-�)�t�H�&"��Y]�:w�k0�c#f=��;�`��j�����/�q#��i�w.w����QS��:�&k5P��(Mb^�H��K��2Jx�����c/S�fdhĖ���!zĖ6���D�cXpK� `�S=�S�h8	���?n#C;��� �n��H;"��id��^Q��N�!��z�2�oL�0t���g�~/�@QTQ���I��T���l`R��-�NM�5A��8��C�J�e��49�Be˴�җ3I�4���.�BA�o��i��D�^� �R8����)A��܀]o�8W�#������Q���E����z��U��X�=Ep��?� �o�����SF�}
��e߫���C�o������ZK#������%��=�E�'����둮�����ܒa2��y�Q�&�Ҏq��TߨfYGgr��t?.Z��V$Y�hi-P��	��{�9`*��;M�p�(��՚3��>��1��l�ǓeK����/�{Az����=�ޤ���F�Sw _Ѕ�C.�B2%~�K��]3��I_��)�Y��k�����r ^ט�N����]�:�<FV�g�Kf�(����O�~}�ν�^!�~�O��۷����u@�����������V*��c��W�⢜ܷ+AuS:�ֶ_z��do�Ѯ
�A�W8j�������ЖCihL�/o7�a5}x�r"B����`�pBLC��A#h�?���`	)��@;/�s-wl����&����b������w���3o��0�'x���z����e��G��!�t���Ygՠ��f �:��rO�[kBe�~���?�m;������0~�~�F��sE�=�n��d�W�����6�Ô�F�M�2墑+v��'�c;�������(Be�����2G�th܆�Yb�����2� ��TQw�l����;��V�f��䓚��
�G@ e{S[#�i�$�g���o��S�~8�����KuD%��C��p�ɋ�m�x��8�ʜ�����*��Y�I�ڛZ�yY���e�d$��0��I@�X�s���O�¬��_�BU��s5	nnh�È�Vr�!�j��_Is[��/u�t��H+�њM&!�bj�6Md��5�-Ҧ�f�+K�$�,IQ<���.��qIW��A&8<u"�������*s\8��U���8��R�K���aKwf�:t��,��˓�U���}�
؁\ZL{��a�����H\"���E��Ym��(�m]I5��;���N��{��f��ܙH�?�s�+�wO%��e�(6&#1�D�.��/�U�2$�j���k6�:��:c�,�:PNc�6�L%�Q���9��������	�tI��l�H��5�]�����M�|��7����Q� J�l��Ug`Ac^��S~�7ޏ`�V�����:NW�ސ��0)�>.�^�k�>Ř��ad�����[z;�4�����(��,Ա"�������Ms��mI���9՟ U��?Q|	�
�?�wȁf�.
�=���1��п�c˝���r��s!liľ�E]oȄµμ�Ic ��]{8�VR	�Qe��d_��$h;^JZR����>&��V;���.�d�M^���]�/T���پX��]�
��ҋ��ÝA��_xtU�2O�y��駛�RlS���wNWo���<�o�a��:�[����\k:�0V$6����ף��쵻�a���6�R��^�����zB��j�s�+�L������5հ�����V|�z�g<L�m�}�g��_>S>qN�y�S��a��m���'��ثX^�F��q]�9;��|���-��6ߥ���]�;���P����0��B��Պ҉��kF��c)_�y��vTA\����L�,���,D��	����W@�u�rL�A��8wF�g1lB�û]��fwv�#Oɩ�{���8*����&_�k�z�
d�܍�$9r�l�s;};(�Ѻ�����6�lc��oŇ��b/Ue��O�D�����殖Uʏ�w� ]-3#��|-�)6'�|Ht�y�q�hQIm���F�<g;���#��w��hE������ٚ��$QQ$�i�8����G&�N*fkv���%P�p���B���:aC��z>��4�XZ�������2�9�#{�-�����Ffǖ�GI�Ǝe/=�EB��>��\˽�����So����S�u�u�U�m��]Y|΢1��JI
�.����ʹ0�����������G��G���B�N
�T^ZN��ԍs+��h1�}-�4�%Ȟ��A��cZ����Y�3j�F���p
6 �������������j�B��8w��d*ޮ��PW�����Șq���gR�fs����\i,̿��#Cx�?�GT,5M��7�(�|���̹q�@W�7�.���S`[~������Ľ�JT���}����ax��D����-��ٶ4�|� Ѵ_3�Y7re�1�J�!+�&lR k�\#��F~�t'�����;���>�I�JZ�)�g$K_g:�cV�)����G��+���l#�*��zq}S�jG|M��C4�_8�A��!�g8��-�̞�T�K����{@������?D����iOy����V<<e|eWM6��� �<�_-���ZT$-dx/�8f�\� ��ǌ���&E ���ʒ�3�ڵWP�~��Y�3��E�|�%�$|;`V=�
pa�"ǳ�)�r�,� �s�AS�]�IÞ8��⋲�i�u΃ �F7!�R,�r:wY�72a|��@[�}��L��t�o�u6� ٷm�������ч+3�m���B��.��Y��OI�"�[� �"t�qa<��H�6{S^G}2' ʂq�sy��`�W�6S�x�q�*S[ɨ��� ��vG)�wM�C)�����Os�ϛ�Xʲ�a��A.��?y�7�Թ/i�A�Ԁ#�a�0$����`Ƥ�"�/`���⮌��&�}�$1Ӷ�-��3n��hR�C��ւ����<	�ޏ�$,��)	uj�A�JA��I����قW�gê�����.uT^�=f�u���c>��d�>Ie�А��j�U5��:`��i��
K1B��J�>���"*���
�_ǒ�x���|��Y[Iȷـ�G_��9Ⱦ����g����,���X�fh�n$���̱�_��c�������7´�i�g�2�#�&�!��1Y{(��Y��4�U�+��q�zq����G��X���n(�;���$� �����PT��q��c\^56�
ot@b��j�۹ltj-`p�'�4�<:�_�����?*�8m��w�ω+z����L�mW�Q��g/��Q�nyv#.Z
�������d��T��\����J�&�'Z���	VJ�����=����+˻�÷�Z���xn(w�����#t]�zԘ�׋{N���{��)(	��	Q�Q���Ll�����=$
��ۖf^�J��å�3�ˉ�?d����gC_�YCX]ǤX{�U�L��3�i�1�R8�G��4�wK�Z��yj>V�;����NA|�!�M�w�$�W�N@{w�����J�|��'��������)bte9hY���'�\���m�y���էB�V�ȡ�a}N4$/��GMl7W�c��[P-�cǬ�4��� 0����V�eӫdn�e�WV��{	gֲ\|��@C�V�NA�P3���cK��F����Nwi2MѲ�w�|��L��]
"�@$V�x)p����xT^:��GD�B�� V��Gtޘ#{��}� �J��������=�3|��"������2W!�J�4���i(�'�8�46����l^��-��ժS�s�\U�{���yN˻7#��P:x�&c�h�p�%j�|Ȩ֕���U�~"r�T���������Z�5q�ڈU��R+.�K3�L���Z\-j�l�V_|MbUXʂ��S��5'��6�ܔ���CNʃq�Ǫ�E� ��f� �+�0����S��������!m��`҈��]@s9��!��
����V%�S�AŮQ�KmcF��ߜz�n�p���Փ�~�~� +�B��H�Q��n��E�.�~�k���E�b�����?�9~��}��p�#�����.=!����/���%��ڍ3��'iS{i�#T��қ�	��0&|�c�w��^U��b�ÜJT  eXG�ϣ�w1�ᜮ���i-�A�3+�(�;�;�m(%[�f��q���ڼR�<����	s�7Vjŷ�:�"�~FxMۧ2�@_?
�*U|S�Q��=w�!!d��Y'�CtnZ^���q=�VnJ�N���닥�]��jT�R��&Ȓޛ�ޫSXReZ��Ȭ�|�U�:0=���`AzÌ�}Ǌ,�h0�edY��i�PE��#�/S#Ù�Y߱F�WQ��a	�H�%,͓I�2	�T��zi����ʦ�J/���V�u+�A�P�&�Vo!=�Zꛛ�TQ{����4(d���CMN$?֡An�w����k�ܙ��`��b�t�.�^��b7�&�T����N {]�b���P1B�Bտ����E����D Q�Ԃ$������烈@�%����O�p�7��mU��F:����"Ec�EZU�ƬJ�hd	M�_�+��-5&�`Fp����^d*�"��I�}0�e&mr�"b�v���z٭� ����ϟy�� �2Q}�T��I����CLބ{���O�͖���is�����(G�S��<N|l����s�G��>���r�p�$s����8a	S��*����-'�Z;�]*�J���s�\�z�NS���y{_���K�׻��Z#Ư-OU5�k�6�{�Lpjoa������ϖ���#�.zV,*�7S#�@�$�n^�j�����vzf�Ua�3aNAS��f~��>��	�����]Q֛_"^ي�>=���iM~A�w�o��p(�{��/y�4�a�&Nn��n��G{5�33�B��A�%)�?�',�Ƨ���M��!j�vv�ߤf�5������^J�&�Mky��sŻ��M+]d]�G�CL�y��pa��y���>�+{;7�l�uMÊ*�����Q����u�W���O$Ʈa����b���i��f&!,)�A�0��b�\�%�L/b���oR��rq%��Q���`=��Z2ᨴo�"��ev[\T�>D�9T��tO��m>aHl�(��U�"lq9%�y{;N��R�k�!|��UqnB���x����*��Ş2�W$X�P#�&��{��Q��w��z{˿ⴛ/h����� �?q���M�~�i��ޟ�����o~ٺ��*0;�/){������.M��A���z	3E�P<i���I��,�:ܔC>��O�1�o��oR�/J�|I�̳�ә�M�q����8� N���W7cmXZ�Y�C�9'���t[0RHp�qXv�'��ւ�8#�TU���{:ԾBx��/��ͧ�o�`���,�1��ja3�]`�Q(�_b�������兡	�{�S�O���f]8OJ1&iw�\�{��)�	�H�?Mq])&�?�Ӽ��&��;5o���u�踯Y���3�.�>�頙+(Q\uDA3�7.K��E
�2����ɦ	oI�C	y1>�A(G����G{AEf�6�����"�z���ą?�vp䣗hڼ^�g�Z|�ǘ�yQ�OG�M�ӻ�o��_�JZ���]'�R��d��P��B>���pjݱ���h�U�k��2��i�<�������WC\������U C��@(���<THV4�
���93�)(��������Vr�Đ茎?u-����Z&�^���ʹ�ڧ�HO$2�)�4ߋD>�&��3��N�E��5!�b��D}���qKQ��8�"�.�b�t�;=7�}�q�[Z����ȉ����slb�YĊ/��M;GuYz%�����;Pph��S0Orjǉ�$�K������?�f��� �u� ɒ%�0d��o��W~�9���O K�K�]����P����)�W�a[~b�R�cs��WO�����8`Cս]�5v��h�$���|�u慴�i	'd}�˝f$ ���Ό�p�O0ڃ���Z-5�X^=�m� �efU��VL��^6��<��]I�BQ<�R"̓o�2Hv2��y>�^;���>~Df����C�����7
it�%�v���K���B��A�5j�GOFY��2�|1�8ė��Bc�"�r�sOڥ�Z��K�G�W��6M��7��mDѣ�a����)P:^M����ժ�f��ͣu��������7�����N<_������pf+�OJN�Pv�X�aQ�	�q
�;��?W���w>4T����.��ī�'+[q I��p�[���:Y�D�6I����}�`ϐ�NsA���}6�p��$�O�֖j	�PC��Y�qf�Ӿ%]ְ:Xu�4�o��B\�Ûm��Լ -���[�C�Q�uï�¢�n&u�����`%�V����*\	�#��6OÊ���CX����']QE��g�W��W|Gq��-���]�9��@��CDG�jM����R��FxP��;����t2�Ư6��%!#ai��O݌�A��S�>a�e'{������PI�Ǵ���?0�����Ӳ(1K7���R~��٘{�?J~��Q	*�0�m��+y���(��h*3�ț�Q*v����m}"�Ht�e������&�j�����6�f����%��r��<8�v�
�s �x '�\�Iz�m���@&\
Wؽ"���A!��X���¶���i.��*.4<�
 ���D	������0��2���x�b˞�\&���_�[�E�Xr�A"+Vx����e��p̂�`�ΔJ����"��`�)��rZ	���% V}MA,	ߍ5x��񆣊��U�l�"�6S]Ih>}ܷ�ˮI���Li����"�z���]��A9*�
)��,K@�p �<���	b��~����)��6,X�KN���fc�$�Y�����!�,�	^��{����(|8��3������k�0�9��N�X�������`�miXcV��17r��~tC�(Xܶ��!�,@Z�����ta���q����mR��h���[��J�x$��<�"�Q/�c��\i�y�u���ɬ�vfq�-��ƯT��R;����H,(�E�,!Qx�܇|Xo/p���ʹ��1�=���9čk�?��3��K�wG	M_�pU8���˾
_���1����9��Z�hF�m�Mx9K��RU��Ӏ9�Y�.����r�@�ˣ٧Fi���K�>�C˵�sp�dY@0�גq��{�f��k. �L~�������^S�?�Q���eL���j��GL�B��i�������d�����6H9L��Yf&�O�6�cUl���/���QhEf�{��U�k39hZC�~\Ռ�ۘ��+V�9�*�]�~K�!�S/�:��h�37�*oAe@Q�.Jm�{���^ H�W�2fLP�@����OP�+���%m�С	�{ �C��Z+�թ�W���]68!�e�I�q��$ڻeH�[$�uĜ�c��hJ���a<�l��ux~:��(?�ƥᏋ��Z׼�l*u|�E9#�;s��M��B/�-��ȋ3o��.ɟŊ<V�����&��%� �{Q
���=�U(�&���g����+���U?���S��hK�����\�pw��9�Ӌ_�l,�j��c����)Ȝ����4��,4d~�7�YM��?<�����LBvF��[Z@@�+��	���@XpYoq)�k�瑜<@���9:��s }aw2tO��ǽr�����Diw��q�#��O��A�b���u��Hޯ~���Gѿe!3��y�}נ�/�1�	)����(ѱ~y����l���qC��{��b�(6��r�ۿ7�}p�]麗;E)��c��LL�Χ.�N�6�
�% "�*/;��NPv:��$V�����ޒ
~�m�2"�&\��b���cET�����{��R^���ն�W5��elK2�Ο�eƺ�I�P�,�o%u<o�0Έ�6�K�����t k%�)/���#��c_xx #�X�	���I�Gy�oX���?�u���(��2`�����7�Z`Kh?²^J�W�p#܌�ܠΫe;�"�uS����r�*��N�5�<�%Z*N�@]��� �-e#[��S�ٵ쀇z*�V�ӒL�f0?@�����8v.s��'��,=�U\D�����s~x��r?�[D�wP�gk�q!��GOZq�<���Aלc|ZȞ`�\�?���Eܺ	���m�F��"quق�Oe�H���cՊd�ך$b������CWYf-[t���? �+��t5�}�Sv�,��� Rٮ��+��kH~��VD�܈G�~���&��XU�nh()k��l&N!Υ�)���d!�f0ct��VY�X�G^�Q)�K���<�3`�Q�s�Uj/�~�������7d�hm��xH���E���o��M�:�?���M�� C/��,��#����y�|ȳ� !<�wVZhp�kM��.���g���w\s��k�DI�I���:+lP󽺈��Z'�M�bv��]ux/d����Y�hX�@�Ι�4bD��+ߨ8�}����^�oW���C�I,�?WX3�ڵ��S�}J�3���h���|��%��K���4�.t�kQ!���r���y^N��]F/���d�"�~w�v���f8�L�\��f �r�~�%�6���Ǎ��inv�U��A}��Mn�t�Ƃ��@7�A�Q��-�9Z�YC�?��ׁ/8��^��?=Z�.�:����s�|�XEu,l_B��l+��<a曝?B�'e�ڐ�wʈ�*��'c�#֑21���e?�c��Y�6,0�����=��m=4t�Ws������L-��ȦbR� /�>#!Fc�)l[�%GMG���[_�-�2��Gt��x}�us�}�ڡ���u�#.L���6�U{�)eI���-,fW��wO�t�4�f���tP~Y��ŋU@��b9dT?�3�9}������VlߑBi
~c�����ջ,A���"�dK���<[��>���]��pn���A�g���zK,/Q[:p4�"��}�:��=k ��F�No3MZ-�W"]���y{ܕxޚ�jD����YBW#��3�,=�����*�%�!��GİW����>�s3�k� ���eTW{��t�Wլ;�:x�Z+"���j����J����Č��`����m(��S��i�D�������%Q;��9pI����M�� Ac����Ɍw�^�q�ܯ �Tq��bw��J�����Ex�D��� A����h��a��r��}��M���E�Ţ���LT�Gx��t_�0����gB�.p�>~���s����y���]�O�q2bޥ�����4��f����Λ�~�U\צ	�l��o���5��`�s D����)\�����?��\�<L�{to�}�f˦��M�4<rO���]Q��=�2������y�d%8�<��]5j�88�aS r�C�o�nf�vf�Dk��k���'$?������9-R���`�7���a��!(�0�sM�)vԹ�+U���<��΀��Ӗ���~c�=��G	�N�dt��
�e�<������eD���}���q�_��A�M�Ա��OԗO�Ȍ�P� �ʧ�D"��c���l���vV����VХ�o��������~�}�%���ƴ�$:��?'+�����W�̓���
7��Q�eM5��~��ƚq*�m�pߴѸ��2{��9@<e�ZxkL�`��;�)'�w�7�i��!s����i�~�y�c�ƨ���8w߰ �6򠢀�ʭ���~�b9B�m�bcx�p�<RcΤ�u��e:Ժ�y�(w�̕z��?8/E�T�s�A* !*�K�Y��5�j|������?U �c 8���D�FƜg�p�FE,������Sc�J��"�����`���C�ܑ�T�y��7|��5=1�9)�3�ʗ��d�*��@ΌI�����n>Zx�
�={bv�B��LH���@c�f��%��@	�\��,jƎ�J��L��b?Q�� �|�.�a�Z��Z�;�h��c$%�ܙu�����x�o��e��y����q��/�D���D��J93�'�_�a{>H��n%u�B㧌o�����8��,V��d���qRd�n:	N_;죷]U�lk[�Hf+����󫰱o�ʵ �oӆ
�ᢕ�p�+��A
� ��S�3r���,�]: ��vaa��;DbU^� �%1��؟zv���� ��,�h\�b�c4u1;�#1uV�C�0�����f��fJV�σZN�P��aJW'yL�pb�dڄx�#�t�c����Շ �Ί���])�j������L��&Gj�+�4�	�4�T�9�1�p�A�>�|�@��(O��H=�*1�;UL�4�{�)~�b�0\�#�H �Z+��Ĳ��k��-¡�ۅO�f�-��j]S ��W0	�p�c����ʄ��0϶�s��Y�\��~L��ps��)~14�9�����K͡)[y����J+63B�}���D����IvZR���!}��������j�~�:�D|�i��UI��4i���������)���`�NZCֶ��-H>�S��I��pXGm��v�=`�����VL�#�!P��V�=���_ pje-�n�,�XS.�`����Sc�O|YFL�x���#_A����<~I0�[�>�x���>�lJ��px��Ể��7�5r�K]��T����fr�6�ޏ�]7�S��d@�ɕ��N��<�;j��p�ō|��ev�����:`*;u��<���~
P�k�'�0��l�xNT��qj���-$I2�=a<N��Zjp/�w۝bQl�u[(�i�W"$ �A��**�2��ʜ$��}����~.���ؕ>C9ĳz�_��$O��
���'�3�����$� ���p�����!haW�2	���x�x���b��TZ*�+��+�
������ ��}���P֗6D���6�  ���o�]��}��#�1t�jk(3�ϧ��(���u�� ��N�8�����&�%�����0��s|��_o�a�3v��Ul,�$ۛ�r��:2��4���Eo��׭��C�
�=FTX9ר$�&O��?%q���9���s�D�z��̂�N�(l��D�G�X�kP��2��'�p�=��~�rK�/�X��`mm�Z�аp
����v�*汰VyXF��'���E����2�TP]��⵰�
F�8�P�����'p�Y�n���gLedy5w�O��"�mIwǫKJ
�5�@wFLZV|��f0��a@ΚJh0V�駞8�{\�W-�ip�~���O�Q�t�w���T�'�S�w.��*]\�B���&�9��]�(>s�Yo�D��ʈ
�Qs�*�B�z�%����s��y�䘴�N���Ҥ�	�⍃��u"`�S���&Ԇ����<��+Hr��y}Sp���_�^%T#���FS"?�j��B�ңj��H���x�_����9�,h�)��(P�Z��`��4����mo�3^�}��D��GT��&��`�0��J>I�my��Nք/d�w��r!��� ���<����'�Io}݃�EQ¬�̄��x+�T���d�Ǆ�/��
.��	�O	?r.s7�
�a!*�������4I���ڰ,�Y�ٕ��C�/:E�j��a^a�xh�b��������G��9��i(e:��_�ut�<<� 0F���)jJ�+	DZ�T�K�h0�H��?(��Ys{����q����`�:�J������­2�������.�r�tT��{�:y)E�06o�L�[�gm�Qp
��qn8�E�X�Q.4i���^ő0R��5A�bɪ��R�˷b8_7���D������r��	�e��?�l�ê����fY�d� q�oy�i������>={grQ~�:�ou�����t�9Z��8a���j�q����P�c��`w��_�Ů*�=vG����/o1|�!�Z��qw�������Lp-])��b<�(*�w�.%:
�4�x)f>��$5>��X6���۲������&�u�}�?���l�I9hg�3�|�����^��dc���|�Ac��t�kЮ��>;�a��ZI�ed��|��zD�v�J��6�Ok*t�d�IŨ��J"�U�q3�*��p7
���3�6�uHt��x�G�X���nu���Dl����.3~��VI�К��%^���kY�;K���5��7� �i*��m�Ĩ�^���-a���2�N����wz�H�Ev�N)���{���r�Ɩ�f��v2�}��B�[���OvHE��Y�����
�s�.�D�k\i�)����j3���-@�\��$��ΉL�%InPg?���~���kH��.z*�6� �|�Dx��ұ�w(�k�Mj�.�z;͏�M�6&(��!n�y|w�m�E:=�Aa��A`�d;C�H@�V�hzX����\+���QSL�b�憈܀eC�~�n��f$�;��l<��i��'���}�3=���MM�11�=R8�g���jQ�٢2��4�kq[���\�&��K R�R��-I���F�_��9������30*��<��;#/ʒ�㰛h%��I�,��4���m���A=����[�6�(���^B��p��9	|�YA�L��,�U����,�k����RH��뭩tv�ؓ3�Q ����Df��!�Xs��X�Am�`�U�-�]_srl=�dx�t�S�~���Q��x��2d�O�71�6�N-/���_k������<!�O�3��I��P	����-�=+��n��G����iL�����/����X�#�
�1=�-@
�<!���z��&��êbd����O���ǆ� ��JGǓ���)N�=�Q����<���Z�)��Z�*(<��Cr��{�E�(�������� A��G=Z�A�Hɠ;!Ī���N(,g�]m�M�M����fhށ|���
Ax��j�rл�&�8/�6�竕B</����쪪��-L�l�C��1�H:����\4n.i$�KS�����详��\�� E��x�pM�!�/�,�=�Pn��&����\!��*�S|��l��q��Q�:%��;����)������{/dxC��,��;��!N�o�n����ÿ7�1=\m��2럪�;�R��I�7�i��I���^e��`�C2�(�t�mi�n(E��N��Z+�9(~�Ĩ��Ԁꞔ�\1ץ/p���v^.���S��/�Y�a�ƻ���M��&=>��?":�����>��UK7������x�V��u/R�����&��"���h�$�Ot�|�ɍF]S�W�}A����� )'R[�CCc�2�o��I1N��[��pЂ=��/2�h�}liX��m�0}S�h)�iV_�rM�Vj�	��7��g���%W{�~�	�[�؍����kmɡ���	�������u��PZb%�Ñ�a�^�GQ%TP���J��j�[���VeT{W�}1�JHp0r�C�9�:��DBu��!u�
u���O��5%�֔kP�$׺��b�^���~W�\=�.}�
�Q�]�t�u��N�u�����y^�\���k�O	�C>V�r7��(���9�t�QFC�Qr��_���ơ�_s������0$��w;�leZ�7����e��;�`
� �K9pZ�҃��1�"�q�!0u�m���`R
�5�a_�P~r��}��/�Y�x6�pP'Y�ma.����WW}N��Q&���h����%����kZ�QWϭ|��̔j�A%�S��!�e��ԃb���=3.��V�E�7��
�M,�	c���C��@� ��Nʅy����d�����s��PM�EW����#�n�rLO�����z� iN�۝x�3dl�T[�����ysԖɑJ*�� .��m7J��޹��5��v�+~^u3,jg)��������ݢQ���8�[���ʦ�y,���fx��@���r��)�z�m>o��*T�i˅#���?�c%�u*�P*&*�-�N�Uv�V,,|w���q�s�B�b���(!��-��]l�7�d^nh٠5$��-�@�;ZW���ݢg|0�0b���E�r�|侸�Cĸ��ĩ%i!Oi#қ:u�v�ұ�ݦ�x�G4*E\|�h�9^J܎�qBʧ�-��P�T+ȸ���D 	��É��N�@�V74�xr:}�'��C�ڪ_��T���!�ii�,��=���}�� E�X�}���9w;�R��(�!�f�@�W�!ڲ������1�$��BLa>�:�'=@�|�h:Z��z�?��cV~�7rTS;���Ţ����&+���\�W$6Em�NK%LX{Fvɩ�x���#0� ��"��L@ׄ[�B������9׺y�]�rJ���̲/5\.N��V�!�U�� �p�E�LdٕjD���	/n%�资0?���1��7w^��N<�PRr����o���XL]wr�xS�;I*���}�L�e���Fg3��A�� ��/�"��C�.Q�O�q�yVbO1|C�YqP��>44�p�t���M�e7��B,$՟�g��Rw�������cL��� ��o�¸�aV�{L�ѵ����R�@2[=gn�B���h�g�v��2AY�"<|Q��z�X�������}�&��|�����m|�w�4�H��B3"bA~2�B��Ty�N��z$��*�٤��@p���(�Tt� z��	�|�~E�L�\l!���9%^��򛄈Rͯ�Bs;_7� �'Sk��m�g(jX��;�k�k�"����f�������}ESz+0T�6Y_���'�	�Tu���� L���ܹ�j����"�e4��V��h鑨��Ⓥ����2��+�UBC*����$�Ij*M�ֈ��j��k ��;Gq*!�(�i���<����H��,��i@kJlv�С$���ªh �úD*�#w"�(-5h��Gn��\5�joXS[55�ir+��3�d:ma����4��`F6FX�{�]�@p�INe�
�6qj���u�Xu����zs�V�T���3�%�:�b�Q!I������ľ��|�JA�t��ů��΂g|��"fT �incc-!%s"i�U3���؀B'i�FD�����`�b�|b�5�h����מ/5�Y��i$	���T�� �M���܌<sg��������rQP3��!7;k��ήv��X�.�����H�5]�A�p�`�_�]eV�������a?!rۯ{���6�q��Qf=ôb}+u�x��<Aٰ�&ɣ�?�b�� �һ���ES�S�@��c~�\�f��}�:��=bo�~Q>h�ʓ����[��?�� ד���B��J�2Rt��R�^�㇒v������Z��$��a,h*����8��ӂ�i�Sד^<�U59y=A������X�џg�ʭt���m�O����] E��FlJ�_��>��%����~\ef�w�Հ�u�
ꍸz�ê&5�(�������/��x�x'\�f�X��a��'�:u��w�^/I��]\wJ��e5�]gZ�L>� ����&������5%�\8l�����JO:��w���m����!
�T���3aCuS��J�f�8i+�&�<���M'�7&N�$���/I#1�(����H�w!�4����20��?؜�@�aĒ�Ib�Q!]v;:�/rw9=��q�Z�_UU����(Қ�vƄ����7M)aV����w��ճ��{�K2|��9�W�H��OkCB !q+�U�`���᝷蛠;(X��4GL��:gH���+�JԳn�*6����oUDT��w��f�p7{Uɫ�u&����f����vn���x��ˀ��;�]`P�RڔS~�e�1��G����94� e��Oo��1#m�������֮yF���v�����T�;)>P� �ÔMwB���#��[d3�$"����%^Ե�!�][��������|�9U��O��8tXC�U�~�0�:o���ѽ����T��nN��q��^�T���8�!:q!��<|>��(F*�"�c���h��A��E�����;/ۆF<�cPa��oQ��u��qn˃B��R�'�X!�`���
ǂ%�A���u#!1��lkc�l��#'�m�A�S+�N�'���n	��T�O\��G���î=�ȡ��k���ە$���!+�z�e���~#`�m+6,�$�`�j(i�����
��Sc���$_9%��<N�p��VZc�/Fq^ou�g�0	Y+�X����(��B�ykR�t��e����$dd0b��3^�f��L1�v�)�96 �f�䚙Fb=,������nPjri\��~��;F<@qow�TԢ���摎�����Q�yLA����beh��������³�R�4�Q�KAQ��|��d�9��S���G����m�� U��:�����,ĩC(m���1H!�M����$�����dN�.���&��5�G�	x���S����Ӱ��k �o	 I�L��!�.��(���XJ�Ł��ڱ8<� �D�w� �����~Eg2_S$�ʙC7<Ʋ�y�#�x�&Z@zD�y^�U�� P��7�50��L� Lm��/(MIFq P|�bX��2��N�H0f��~_�����qH#�!��i=[gXf󚜝�6FXq�/��� ��A��W���]<p���d�8E:��]: �o����?�80��_|��f�3�I+���H�.%��:�X��[�MV�C���Ԑ�Y�M?`�s�t�[��{'*��,���U/�$��yK-��Y�f�7�@�#�����71�Q����!n4&�Z�9.���3:XC>��G�:|�|��<x}UF��'g�	���4T8�#�-��w�rل"�>q�JV�wpW�f�`�^���TA�t�N��|��q�w�J��L�?%�#���u��\��~�0R����ؓq��7q�#7$�ν	���M�S=S��a%@#?Bpo�+�*���Y���^~÷����d��S��������*�>*[��R���y-5��L2�+��$F�����d��I�܍�M�#������x%�i�B��ʐ�vGQ�޲��x�J�%
�p�F`ל��%�
��Uc��&�5�4*5��Fg���!�'3c����y�����w�z�W��|H����R���!�j�
�� �)ն��"�[�ȣde�=f:�s�_G椢�j����Ͽ�\8�����[Ȧxr��c+���^�ٯ]��[z�f����_q[	��gO��n�_ʝs]m(��g�]�g�)�`��5	q)%ג��K��@�nh��
���R�taC��r��b�I�Z�I"��qo/i>��9�W�?}������\�;���?7	��MlH霣� �I�=�ꍴ���'��=ʰ~�A�����٢~��8���P��OY��K���J���[v��[ �xo�� ��4El85z��z��:"7uo�;�S�Kpm�zUr�5u�������$yӕ��x���=\�����V�T��d�LoTw�����F��-}�nT�θ<6$Q�*��9��ݱ�H_�)>Pi=�y$�R ��"����ޥp�.D��im����G�a`�f�� ��<��J�8heM��T�4V�'��  �X>�j���4��"<ZB~H��H]��#"���[_���\`4��C/q�X4���ϚC�'R�";���l%�� ��[ܘ��Ѳ�	��%�Sj���V���7b&�j��7�N�ߺ�[��u�CY��y�zn*X6����jf�D���ЬX�?�Q�H�LI�na=5#:�.��.���{���1�5\�Η�/ ��. ��	%g��6���^��sᢓMR��@fG��+J���['S�=c�x�L�jO6:I�k����L��ʵI���9����mO�Z��w�����i�����y��5�̻"47P��B�(�����r*�q������\>���5m���-�}dnM����DPT������S+��.��w�u�E��|�2���S{�hN_�H'V��͗�Z�ٚ�7��S){y眬"`Y����>�j~ˎfܒ����\�����&X�M�+U����C����.���	����ם��xUΫ�Ut�ԑ�[��p]��VfM��(Ӣ3�N}�h�	�]@YO�H2�0�V�Ǿ�Д3�ၾ��sƦ��5VK}���+��۾ң����O�,{�Aw�!6ƾܮ��e�k��b��xc`�0�'-h��H�c����.8����u=[�������aj�=ƙM����pn^c�Q���Y���5礖�I�L�n<a�90/e��-U����r�N��s��b��r'�6�z"���I�՞��1�G3,�c�"��T��M��o��$8!��akK�q�vo^4T��]��uۀn��$�Il�g��;I<��S4�}���,;��//�g��_�]�,��_0f�A�3X䳾J��6�G<P�� �I����E}+j�����D�1���TάY|�=oÕQ��I8�6��x���z/k/��JW8��.��2�t�Lj1���N��Ԩ��Mis<q�O�bؗbO.�**��dkښl��{|����w��0���"�Y'�6�-!=xܮlgZ}�� k���>ۇ-�@<�~&��V�"���i6�aE�q�#0q�����x�d_/M�tW�lzp.����^i���0:ETMu˷�ґY^�?Z$i��"�Ȥ�%%:�\@o[��t"���!S\w�|Rns�ٻ�T��0BJ�,p]�@!|J�&�x�q��i���bN?;:I��^x���ڃ�a�22�wx�D�],�V?a��CC��{ԋ�FL	���	�f�:m�"/�Ocn��ϴ�;���T���C̈���|�%��m�bs�J!V3�$GcF1J�Xo�ﴦ�>��}_˼��V<�+�������*T�Uv�������0�S��J5��vz0��(��l�Q�i�hdyc>�f��n� [�J t�#�Fg�9��ލ^i��/h��5��� <�4`<a�Vj�2z	m��~��B��jQ�F��B���g�����K�U�'2`*V66[���{PI\��n*�,�]��%A��~�a��v�>���"w�����<4� �=g��`�7��lS|����d)F�SU��?V�'%2�>�"m��b���?]����X%X{�+np��!���0'~�<�\æ�m��� P,�n��7�5���l m󉼫.��>�B�"gcӗ�<G�5�ז�-�w�S���n�ƌ$q������D�̀�N���l��P��-���Hc!o\�w˅���z܂���V�cS��C*����sG�/P^��װz�RN�#'����ї�,��iO���|Q)��9���7m������x�M�_�S�7P
E�P�*&�&����e
W�+�謷
}�%���Ȓ}�hS�$���C���w"��M���
��ΘR#w�*�c��;�AᏂ;;�.j����Uh�X� ��$�
2�.!�A��x"CHV�"t���v�q�������{2��l��MX����h�Bt$*P���	�9g���<,� _
 ����<L��d��q�蛴�� �eD�Sa�qt3�<F�/2�br;G2���� ��^$���+��VG�P��x¹FT���ڙx������
�����b~�>Ԋ�H��e��p�{��V1���]���o��Uf����K�R�(�g���Nz�S�"���<�:G��ȷ�;ܕPb��"�� ���]�q\���_��/��_(I�b��'#k�W��ӻܡ��Kn��O�A10������k�)�j�y3gO�)�B�_5^�/ncVX��@���_:`WF�q��c
T�v�5��q�&?2�Q݈	?�-sn��Wm�G�3�ֺn�m�����"%cɣ��'��mGb<ݴ̍���ӏ2v�i�9U(���0.�FjyN�Go��[-�#'��a��ǒC���Me���>�B�a��b3�ݨ�k<8w�j��� (�����<�O�KT�m$��Fz�M���빇Ic�,&���4=
z��B����^�ֱl�D�t�9��O��(M6��1W�?&
pS׬�T1)	[�ْ��}~ّ$�G�pš��Ơ��������2�6��!ǜ#R��;�+��7�#PUs�͖�����D.1+�N����ۻ�I͡#~�Ϋ�R0��gn�y�I;��ƒ} �V�%Y����8HB�`�����H��oAE3ʸ�ce1��o���'�Y�V��T�L��Π��^HZa�܄m|�^��ɻ�.�Y��q�b�����4�Mx-
i�R��`�A5���;�Z=i��n��W�,W���8N��ܔ+D�:f�H�5�B����-z@�.���\vD����'/�<���~���'��[�����6]�]�r�'�d�R��dp��jeh�g�VAk��"˩=ސx�+�1�Vѣ��M+ȱ�'�M�+�8 C�oB:'�k���hd�\ ;Akk6L������d�p����섳�*�h'7�gh��ؽzF�K�vt+n/�װP�qN\ҏ��V�vG�m$$�t��KD�}m]%�m����2|����K��Y����Y�X[IU��y4������^�!�Z�VG���S���tG|m����<�j9�~�/a%R�۝p�ag����R����z�BFFi`�fk0n�2K(@!?\�r~���[�&�s�ѦJA��a���l�t�.8=�Bm���;���e���o�A"��l; k�4��ۘ�$4��tz��I�eizG ����<t�.]�q�;���D�o��%�|�Dp:lc���CL2�'6�KV�ӪQ~��� 8)5_(��wL�c�MӉf��EOײ�wW�����>ih&��bcA��k
�S�!a,A��o$i�3g�׌�	��D,��W�)�������'�х�,t/�����&�pbO[d��a�5��$�к��B�DYI�[bv�q0�r�_ՕBF��^�&
���y���,��1��ʂ�)�+��p�B*�B�:g��]8c�Y��8�@�k4�I|��1���"�I{w-��舏F�֍顈Oś[�0���b��Nw���E�\�:M[rP!I�b�g��-���?��D�SZjF��99�u���1KI��Fz^��Y�� `�)���E�!�k)�	i�v/Y'FzF�-e�B���)\y��͌�W�(V�t��_;dJ*�(EC��W����:����\���#�f�]�4�l�=�`� SI5/=𼸱�������a��)��#�x���r�X[� �@�@[J��O�y���T�>���&�.���r[�{���+�e��<TR^o�{� LH�/7��bj��K4�[a`J�a�9���*=d�!)ϹY�d\[Z�&���@��K%|�p��}�a�T�l�y,E�[eNS�,����8�T��sX'�I�^�D�Ѽ����c�2Ism�?Ӣ�-����A���Pծ{��cS�L�!�޾�T!F�'���`�}/Y��]��']Q��Ꚉ����¦h�s����
S�ʴ&�?�.w��Đ�򠢾�5��8�KK�n��>a(�6�Su��V�t�?���ť5� p(J7����Yx	�}����#��g�HJԽ�y�=㜉�._-8��%Q.���m6��#",ܨ�#\��`1{d�VшS��ڕBH�4��G�r�r�\r���M3��4��')W�B��Y�(;��!V�祳Ժ��vP���o�4����Ulϲ?�R�|�.�b�@v�P�+�D���5'�wG�m6��q!�*&����a�єk�̨9$��$ln�H`��<��������]"��R���ճ{ �a��!��obn�͑ܞL�ϑ6��t��0���6K;�ci��bzsl���v�^��~H�6!����4����l��@?�`j�I��S��@f���M��<�A6 7����Ȋ5�)]Wb�ґw�Hi�E�P���<�������kO�+�)�T��i�I�ج&b>9�٫}��6�bDU��N\�Q���gu)dۓ��a�#1:I��+��0i�WlO�l[��P[�E/�}������=
C��sx.�D�w��T:]e=+��:i�:�݊p�KMi��W�n�YI�T������X~�4��3�H�~�A-���EP������"�'<W�툕�I�g���fS����Rw�2!e�A��'M���������;0ٶ8!���%ʵ�O%����}�WQG ���o�U�D*�tө�[h�	Mc"�zr�^�;�[[�ybY~�O���-O���w�۷b�O����%{*�@����5�h���p�e7�Y�5�,���c6��9�k稱��]w,I��#��V7%�������jE�j� N���c�q�<�0�D��@�)׭0�2�PѤ��	|3�_��d�Y]�Y ����Z�@OV��kJ���uyeHn��&����E&`����7�my�\dm�N�5ž�v}k��͍�uqH2z�w�:��ة�UH� ����?)k����v�N�ۣ8�D�Ǟ�5��3�L�ӊ���-�0�d����S�*� t�����E����41�Rw߅�o쾁�Lh�$��C��c��D��m�RS��i�̲�`~x���+N�ĺ��}W��׭�h-����V�����E��>�ȂAz���eh)w�3�����ja]��%�Es�#k�E`E��`*�Ԙ�Z�&���p#@3��5��K�M�m�}b���F1�NX�gw����TL�x�x	��X)���TB~J֦����P_͊�~�$λ��$�4�Rme��"�nR�[m���C���J���};*�*�lm#�4����i��x��w�1�g����?%���?�E2-�j8���õ{��<�ߔ�ڭ81��nE�4�W�=09��(��j����8��/�,�~�}���r+�m#:��Ar@��Վ����hh��.-���n�V��C�ʽ.�_�y!�\H�1�֧������MC��r��v�:wN����N��*̹H!<�k@��g�ض^v#"�^)���иJ��s"1P��w�G�(+��@οJ�28�)�'cK*��u���x�ܭF���h�u�Z!��z.E���HD�F�W-���r	��5N���	f3h���K�E;� T��	E��$���Q<gЇ(3�7g��nNR�^[��Hm�J���Ɓ OG*�����ÌPN��r'L�%�<y�q��(��܃��O�R��5�z%l��}�S	�~J!·����(+�}�m�'��|z���0��\	>mX�딵��uY�T�B�5U�H3j��<?ǔ�T��a���_6vU�� ���:������Pʩ��5y7�r,!��w�/�zn�8��C\�.��v�i�ɨ�MW�ez���F]m9��Q;�Vn2���h5(N��x��z�*R�U���E��#�B�(:��^C��
���W�팓7�W�} �,]8���#>Kk�_���(]A��d�E��G�'rB]�>ᷬX$7�Bu����Z�������Z�g=w�9�[�.'÷Q�)�u��<*�>]HP<"�L@�$tON��^>�}zQ��|��N���@N��!�H�	��j�;4|̞ڀQ���m4y�C>�i�����
��ˎ�p��!��.]�c�V�3��T<�P��xU�R�:�5a�m��~��E���>��I���9ؑV�d^���!�x:ON`�ԩcx�q��݈w����<!����c�W��#i^��ϫ��K�%Hک:H��&8������L9�II[�yRI�~;M���A�{4fe�M�4M {�.o*�lk���4�ȝ��]+Jq��;a����h◷�X��J%�!�����c���H��v�2"N1��O�ۃRJ��i�=^��6B$+[]�u�eH����+3F2�V��G�T�t<O��]W[5�p'��BxA-��^0�7җ}�)V�'���^#�A,P���4C��U���`�0/S^��Z��:"�vFZ�#3WG�*���^.9 A|�ٍTt���������侒�S���=E�?qɮ�D��q�y�Ϭ��P�n�t�gH�_�I��R_!|\4��K��8�2NUH�5�K~M4��R
ٹm��C�/
�A�j�"hy쓴MVD���1])��2h~}*�>�'�$Ď.�q�f���z\����	��m�5��J�t	N8���$^�{�U�����`���q�4�aR$�%�F%E}~�+d}��|���`G�1�rvP�	��&�����O
�z,�G<��^������C�d�0T�O�Pe�֬�M���O�C9	~�u����E[.X������}�D)�/Q�;ev쎣ߩ���)9�0��h5��}࠶2E�ed�p���\�-0���l�r6�rj@���E�:���a�d�.��#Za%m�:/�	�w,�u&�襏���?��/��P*�8q���a��Eu�#���@4�t��P����	��4�k�cnd�H@�۸�m�_��s��HY;Hvv 
(��Z�X�������g2^b���:
�T3yЀ?���.�n�4n���E�†�aU��WH���]�vK,�0Q!�����XY��������L����P������
�jv]<Y�k�~�Z��%0	��~�E��4]������߯Ye�P��l8��f��iCBzj�Sj��)�#ƫ)�ME����,�Ŭ�׀��_���y[ş?ɩ1��U������6aL~��:�a*^�6�,������SPY|p�I����N�L���`5~�2R�^T8��16m�DmJ4���Yx42�f��K�S�w��Z�[�ף�[���l���tz�`�8x�:����"B�n*���M@b"f�+)�Е>��
�8C�l�C�f�^����1JA;�,s@X
�<�ӹom�q[1|�+I�.O5�7W���%����
4�V�zT��e����"��s���/�o�4�O�Ո�x�����I&�&c�3,���k��فeK���O����V�e&}躗2^�n;��߽���M�T��n�Uc���mif�K���W�g��l����)_n
�H�����}J�_������h�ġH�2g�p��}��C��1���>�����N~��%�Ku� 2d\�&
ۢ����坎�$� (��F��k��N!�����f'V�a��|1Y�x_>g9���IO���t8�=>��)!z�	��%�۸�n��P,�%���Eۦp�*�=K9����6�g��O�M��R���
�J�y#��K&�!<�X�4�9.�̐��F��]c�D��A<�}��y
 NSr;�߶]:�|�Q��z�������ёY�_G�������5����[]m�St��-&
l��@^c|�$J6�H�ǰ��)+1d�m9-�:�z
%Q��Ό�[=w�5"���]�{�J���j�9����}щ�(�(sz���r�g:������V%�껲�9� ׿~'��L�Y��[�D-�,~��ڣ�,b3����T,$�/�R�FQ kp�%�[b�� ���}%܋a���D]�]�/��]h8�n$���ӟ���m�`[; ��#�y� vO��D���G��4T�x���w�B��⏰ab�"��ЭX��S^LfU�i�E�B�*��2@�nc�bf���\
Ý���%#L�м�Ҫ�\����4�������2��*�ϳ��-�q���[A)+�����T*0O�o:^����kj�B��w����\��|�nS:�nu��m6���ݧ��[H��jד�M[;�R�$R9<���.�B�m�/����mö��۱�z��>�꜅������-@{,����+�+�J���_������Ky@T�t�7�^�3��|�ɜhK~����.K��;����p�|J���^���1�oم&���U���n����e�e�bY;X^�!LR����	��qFKT�=�H5�J�T��o���0
W�5'��:,MP�0��B���w	ȸ�����'m��>y?���͢Duü�Q��u/3
�إ"֐!C�?��v���8y#f�i J� S{6)'I%����oDnfe��Y��z9��j=�+�A��rM��K�ᏳI���H'�"�>A4W��5�i\i��u�&e��c<�q�Q�
+�q)e~���Lr�Z-{���	����+�Q8#�ތ῵?���$2NBM��b��yo�	�t�i�S��p�D6��t�<C$����b�qFT7��;>�����۲�^�N��i�q��X���������{���8w���Ic�/�*���;Ri��x��y������5�d��F�$F�Z��y�?r�)��!n���6߾���K�*x���� t�����z���x=S�w�ri��)�I�|��>�wPZ�>�X��+� � ��J��m첫N������~sk�Y�[I>��%y>��	�-�P��%i�,���8�G��;��'㺦�96v���f5-+�"��<g5��m�
�v����t�ɳ�B�A�.{�����y��<�I�8��7��Q��\�5m�
]#uk�q@�B��'�^�LCt�j�Q�d�AQ��"�Go��(3��-�ތI��!U��5^��Z���0MX����S��c������j3�l��+t1�4@\�o��?�\N�?����%�@�����3HGע�ɿc
��4|F��(,,ɺp�Qy|�>�z�尿���NSN
l�5?s��-�O��nz�_�zs�~���S�ϊs�4Hozf��w���@5W�k�դӽ��nNx�bI�ګU��׾�$ �~�M��Q�T8 ����'�g�� �?�0��k����1շD��:FB�$L*�J&|���f��\�T�ΫOֺ��16I�e�`"�d�����A�A*Z���D�a�	�Z�\$���I���lʤ����6���.d����m\*.a)���"P�F1�o@�1��CX��(G��顋�(���x����X�
�@-9}�y%�l=�����48�w�Wŝa��)�`�e������1�'@�-�)����x[eb�s�#n��G���Ѥq���V%������F{�P���0�+���@�f��ӏ̤���RO��/f�Ю��|n��H7�㷮��N��U�G˶�A��E���A��_ho�~��onA ��2�ێ���e�OG5�;���n�)������d��t}D�ː|�d�d�
���y��ڢ.h*�H;�t���2����P�_���F�*d�U�qI�8�K�{P���%ft���� ڴ*<�8��:�ƣ��d��L���R�݈V�X�@@����up���n��k�m_#%���چ�,��L^,Jh�W�aV�:�.�|�:ĺӠ�"y�i�L��݋��Nh�����| �	.�r�K�1ސ�0Y���~��dީBw��5n�����M���ʈ
�|���m[G�?����n5����/prL���`��|	��`�ʷ/)�v�:�;�yѕ/�O5���^��J��v�DW��H��s�8�N�&�8��@l�0������!;)�?��8�/�q)�3ŝK������:ErʸG�	������l�Hh�>���Ǜ�����Q����ߞ7�)/����R����qG�S�Ց]d�|(��?XX�;��AEU\�$v�o[|�`�":Xw柎΀�B�Z�f���p?�"}�uh��<G9����;N'�&5�R*(�T�@B\ޱ���N�,�w�]�^'g,G����}�w�|�|/l��Z��"jo�}-
Rs�T�������^��,�D)r�:���h��V�.'�tI�-�F�V��0^Us�p��C��0������6�35�lJ���������q��`.�}�e���Da�ahg��j����,��;׾4EJI�x��)��م�ݝ�eċKp�da&�&�6�Y����!7(�J��r<���J��L����E��
�����qG:مJC�pRŔ���}vV�N���J�\c���%FCT�c,�g���k�����Ƨ	���r��%N��)wA����43#!��׉�#}x�����x�����@�c�w$l��`��`友��z�Uw\
n��]�e��C���*��;��4�]�L�5:����j֫��E>��ݙE%ny?�r�@h Wδ��\����R`��Ai8�黤�D?���4uM������IZ�/?d%;�N��F�6������H���/d�*)��ֈ �S����6H]�d��+��_�5��|��	I�����8G���Sx�&��r�*��t�������L�~q������:��j݇� {�fd�pbbKV����Ҭ[1C�@�r�#\�V�OK�Qe�ٷ��R�Q�H�[L-`�E�|�ATB���v(���OM�*��s�:��gC:q�S`h9���܊,��軰&1��f�C.vկ����|��?�% �mq�[ ޔ*L#�ъ#79��XMr�E`�e-��s�����Y8s�OGS!��kD���*��Ƭr6�0~)P=>�vfV8AE����;�N��G�H~q���\r@�kȴZV��4e�F��0�vݖ�5�TʰإŪ��<;�!��%^̑���f��E�]��PyYq�}�������3L�޵��!�ԇ��Z/��z��I��<�7��h��/ 55,�0�0���3G��5k�ǎ`w��Ee����3C�겾aR露��$V��k���'Q���r4�Sn��Uu��F��RT�U�Ln�P՟{�)#Ց����.��q�X�{��Y�q�4��$
%	ʺ)-M1W�h1�:{��,79�ENo>)#�
���O�X�z���J���%(fE���ؚֻEU��=�olS��N���s��s�H��TH�k���W�4X�!f�³Vj5`9�MX�'L��?���B�@\� ��5��V,��N�K�{�4W��<#j͜��6X�ҷ��jL��#j��Ǣp�z�p8h�8���cg=���»vD�,�zz�峕�B�c#Պ�G�n'���=Z��#��DЂ�)����D3;BK�%#)�����#��]�b����ɃH�˂[��>�0�Y��׎��U���#�P{i�k�Q���'2�ѭZ$��������a�r�C1�u0�5��%�}_���5�;A�!�ܽ�0�v�t21�~��^��=e��M�q��X�O8����3��n��Q���I1��b��_HBޢ�\ѧ�h�����m]+<�y���1)��{�W^��Vw�"C5�����\Hx����p��u��f�D���)��K�7�ѥ�Q80�p�`�J\�P�\D�/��L��2&0�<ێ��:^���@���1�~�떡``�m���h،A������s��6�t�1�]�C�J�>�qǧ��%xyұ��+����(�i�V�=����.����%h�������KT�3��&��*�2���5U�Gd���ڮTb#���N4���t2�h��	�@��A	���{˂4�Uor�����"������ķ�ƶ��D����!��-|ըUUf�¢��˴ $ܛ��H_KȆkm��_�v��O�����Գ�!gM�G^��|5^�)�Gחk"�w�mv��@������0��0�n��Q"�~B��愰Q���5���ꓛ�.�R!�Q-֚(�'����
�w�:��w��րl�P)���3�(�?T/��#w��d����d+;�uM��_u�
���4&��������7�s���`=�:�Fy��>�ۃ.A�L0B����O���:+?Eq�zT�ku@��L��tt�=#δ���{'"�XI⭋˷�1R$@��qz������R���g�����'���ϙc���~��Ͼ�@�б0 O���+PH��$�;�)N| %z�&�B��R�ݍm}�dEW�/oͷR#�/�a������9�J�F㐃�\�N�=�>ҋ.�52?Q�+_�X�)ag�_��$߱4����G��WF��i�?l��׀w��D��c6>r;&��
�屟���!��b��H�����G�(5�<vvaS���k1�Mj������h{��¬)��~0F���VwJ9�
�i��u\wΩ�$�T�Nxn2}DP��2}�-g;���oys��������a؝�s�@���$�Ĺ{\��o�.�������Tv�F.�bq���X֤�{��2j�Թ�LLx�̼�I�������2�'�l��<�#�h��q	��wsL>gY4��um�+�#劬�B�i���tD�t�Ę�K3�mAZ;)Q�� �b���j��;�$�pV��2�kSM�;��X�i�R� U��?�"���:E�ޛ#���m����r�C�� �� �SO�⍵�;Z�V�<��@��[Z ,��"�N��帙��E=��`d����OI��XLܽ��@��ueA��A���Cs}�I��O�n]3�~�(0[a;̜2cۓ0���������q}�f���M1�����EzK�}
3J��'d��$o��ndE��FaUBh�,�2��M���"��D���7v� AM�X}-|����}�G�_:=��́3\��9h�o~����-�іV��)���%��%���X��-��M%��N�����WM�%H�'�y���m��M�8�D��چGi��/�2a�����%@��_�-���'���Yt�W$�m�;H�˥CyZb��_J���
=�TP�F���}鹷j2`�Yn��w�fn�m���CRB_Ͳn����� Կ���c����8T�GA�������s���6&�E��l7��8w�^m���c����RGDԟ��od;�&��$�V��Nq��߫��՜��_�x�4sUf����g-�'�l�EӨ"��B�'��pg	iտ���j�˚�{�N�/|�W!��j}�������)=ۤDh�e.'�i��s*�r� KC:G'�'*F;���N�'�bq���*MG�z�0���î�?e�3�0Zm3Y�p�45I�Y�����Tզ[2	r�;�ٺ/��,G�X9�L����s�w��]4"tX_�$��/�s���|�~�]�YJٟpE_�{T�PT"q+n/ڠX�!��]!w���ֻh�F�S��d!���`j�Jrq�@���{�����1L����O�RR������R�����p�E����H�k�y�'nȘ�$��94 V:���T$F�k��F�wt��eR_z*��+�3Xk����N�UlYA3��$(��f�'�ߣ���̓����փ��`(i����lC��`W|-ґ���Y����r���R��L�%����ט8��L�&�I���'�oZ��Iu<�	�7|���7f�2#�N�|�kJ��-}ED|�����K��)�����#{��%�%�l��g/���8��}��Y>	�^u�e��^��+�����j$@No��oN��s^߼v�>5H�)�-�>���'v<�b�Jܸ�ƒ7��a�|3_T+�s��w���J�Q�����O�u�7�O(7���+��P��ь���ߓR$s�������Y�Q��S߶{>j�����C��û�·g�0���eP�x�F	����A��Y`���T�J����������Z�=04OЖ���6�I$���n��CX "��~�|����!'d�&P5�,�Y}/
f�M��]��x�D�\9�|uC���qʿ[Ѳ�"���K��k�xaV#aKu*��Zh������m��nA�VK���1c�O�L����y�2�Ɛ���&�`pd�k&f�M��� 9��ג!={�6��m��q* v*�,c�rܾ����
�z���x�J����ִ���m���6��"���m�c�)���~^2�d���D"R¡���3zT���,y3�e����.�&1L��\�DoS�i�6d��?,�:��ICSF긧SM�ִ;}8�sT&��DX$~OgpcYy��~g�� �32��Y(�4V���c�O�^�*B�t$Q�]?�Q��ըR��p��0v����Z9�-�!�E6�JO��=t��b����5N�
�B�M�I�$if��q	���Ѡ����h�uF�q�ևC�a�yV*0��(���YH�>�@T��j�t�XA��Ge���x�z%?PI(����T���li)-�|������M�������=lgHT/�|��wy,�Di�ZA�
�J=@�c�j��h	�M���B���#�\��<V�9zS�ZnŁ��c�'�p$�?h��Eb�y.�@�w�N��(��ő�K:I��6{��S�:�͢c�y�iv/��s�f$e�:�}`����{�ҁ�GV�2�;u��5�*X��g�1)Z/MO��9�L�Y{4���L�����4��{��:n�z�8�8N�u��]b`
�p&5ݪ�Pu��k]44��NZm��T.i��\���7o����Y^��%�&�/��+O����ev��a�$�=-�)�5i����}� "qW���B�+L�yY�4[eSvBAG����]Eр,X}�`��F������^N/���)��j��\�J�'5�#db3�c̦b%��yH�G����T�B���h��@�ؠ��D�.�_A���MU���O(�K��⩒��-GB!϶�A�~l���*�Q��Q��y�R���;+��ω�-��,}��`$A|5ķ1Um���[�|$��Sv��'��Z�]��n#ߌ�P�c����\��֠�[�R��8��UX�K�f7�6h&u��u�Ͳa��V�3%��.�1����z�U�\����T����(����=,�(�5hQ�PP��qoj�Y�����[d�42��ǔ�Z�?�}HK3aL+c>���q%/k�����h	J^���	��R���'��(<�� ��M��;��F���Z��\����sY7c�0Z��f���6��o�~mHRɲ ��;c��J�{!B�xo�H����gs�/(�D��
����� '�G�tW�=5��O�:�*�.�ͻ�~�WG�#�%a������%��C�[~ƌ3�uu5HVq0�x����*`�#��@_e�!��%��
�K΀��#�}HćnЍ�A
3&�c�E�F�.�]�h�Ⱦx�/ܵ��(b�eɚ���(�e���-!�3ñ��!�	�B����M1��m6�W�2G��;�2�`�� I�
ݭG�yww]���+o��0r���7�Eú�JZY�S�z�L�HZU��c�u�u�!Kl��f�e4�B����,їe�Ty&)p*ldJJi0�BR�H��!;�����G�7�m�$�
�ԏ�H��6\��%���5戣l<�"�9*�Vu;��S�W�.W�Jv�q��ZK^[�qA�j:�+�GHl�=��zQ����D��$���;��E�م6�`�KTٗ�b�s����.�t&�aW�(۟5;���.�Ftv�z����q�u*� J z�'?d��X��j� �aO�D|0Z����u�?�O�7�;��q
f]��������I�W(z�Ň| �}�/C��_�����.�N �J4�
����ۢ�za��f1��O�}%��ݎ��w�#&,��Kv��L7��X�_-�=�?@e�͚v���s0�
��H{�`��HC��r�Z
�'��?�Ŭn�m�%��M�� �#3h��Ny���W�bo���Nt�C�4�K7�J�s�+`����T�v�C�ԟ�>0���@�YSՄ�����Wv3R���4� ��6��O�q+'�����ք��!4�IaG��hSZ\�_!.S*G�Ҋ� �������k>&�1�YT<�4N�a�_��m��!���j��"��'��9ĥ�����7���Y7NK.�+(<+Fª�\SwN�J��2H�O����-~m$���	e�r�,��a'�+nax�y�1�c=�)��j/.�\��$o �1�C�ۨnf�/�|�?_��_�&��I�!��L����q�	^�����y�r;g�DI���r6�l�[��p'�Ic�'pH뻓j�$&�F�vZ�L ��7r�jP���� ��<F��gT��u�v��5���w� K�}�b�9��Pb��i�	p��)����I*�*�0а{d!rG�M�T�bZ�`d�1@=�_FHFB4��1kN��~o�`����ˌ�s��p�'���!�n)S<�YT��\Ԕ�^C�b���0��_���W>�D�D���0���@
��9�
��v6���f��&����(�����-s�zE�]?5��oB*~�0 y�_]�?�h{�$�Ge�䳈��4&��~���0���r�w���#�|gvin��XM\�."���LA���/��('O��V�k��Nl�%<��#ߑ�D?-��0�X����+�=-�0��&o� [a/ps��9��6�Ma Jcj~�ޜl���&������ld���.�n��=6 ZU9^�pSy� LFY�e�A�W���bQ����(HJ!��#��e�����/�i�+���$�̖ן"�Zp��F'PL�+��&"uH��ve�|
��P�M�2���ڝB��C��E��|�h;Y݌�-39��#��-g]r�i,0D�M(�lѝ�9�p^���}�b�F�t+�R bo���˵���e"(�<�2����?n�W��������Fd���A��x��4�fΣhY7�YI�����!7A��k�[&-�"��q.ߕ ��Z����J��Y<S�J��d�Obe��:��<f]����T�-�X�.�5$)@g��1RUƺ
vUW��s�(���" 5���cT��G�i����P����ݳ���S,UI�&��2OlR�����a�;/|���X��\���w���B��$��Y���ҝ�g^%#R����Y�_	�Is��yQ�jm;Z��ў���7Ha���U�fRK�1.yL�eNu�\��
��c<�9���7$���[�C�,*�K����LIb�k��4��LtNW��ZM������d���Au#�F����,���چ�Zՙ	�h����ה�`r�}� Z�������-1`�s�� 3F�x]�:i�*�sCv�J�%Wz���O��u�L#tg�R`�D>ہe��"��fЍ�Ԣ1Ko�|�~�����<����Ѿ�A���FOL��(Y^���M5^�A��L��%.q�����/�d�4?gH�fN�8�g��������(���g_8�-��`��;o��(����k0߯�����%�`��b�B'�o���?zOފ�=����L�53bߑ��;.�{��9�B�
����O%��TQ+W�Ҧw�B�\o�_���38y��(.|T�`�w�BX��1(G����F�2_Q%Ҋu����Q���M!6�W��ef�6}�L�Č���ﴙa��Fh�c��'���ػ(�wx��&����Pq�q����s�0l/�0� ����2��R.��o�!�f_��	cNi`&=F{`���,�c����2)t�R�0l�Q�y����N����
S��18�\WH{�Uל?�r��4��}������U�`�E�Q/)cȋ��C�L􋏉͗w�7�n�a�XR'�د�v%�C��n��rE?@���ͷi7'DN��'l1�TC�ar;�Rr�$��N-���U@^b~�����=[��<B�I��>]*��ߣ3�M{,���%��I>l~5���%�0�E��p��7�]"m
5Yp��j	�ouy8��-2�x��Mx�1u珱����,���wd�-�����;���{�X݈���CV#����D�~ �c���L�
n�g�,�{��Ma1kZ�]b�������_�#�<�M�x�v�<�j���B.v��ChS�C�� ��x,�l���Q���*��ac���C	����Q��h�������n�4-ێ�qy[́�d���ר�P�g�Q0��H�'��.�BS����*�� 4P��l���Ɍ�]3�4�[Z���7��_����w�E���WU/�K1.�Ӿ��J�;}��K�l������ܡԷ3!��	u߯���ᔶ�#��뎋g;�Y<1�{s��A��F�c��$��~��i0���N���]�s�Pc���D~�ϛPy����+4��f�����"l��A~�;_�#B'¾ɳ"ƛ �F�E��"\�=�J.5��o���h�On�=�Q�n�V.V�0�޵�kW��1��E5�#V�������p}��c%6��r�$T��v���ee&����v-c-���AN)���yJe��V��^I�ӆ�W�)�K��`�B~��a�� �>B�)��}d�eA��8|��6�&�v��	է����ٻ����˲�)}=J�k�W	��c�Tꗥ^V�dZ��)R�ǚt1����9�hW���a�.��s�As���� ���b p$y�u �/a��_��t�@��#+���Y��X�~�`��-<��8|��5�Ei�Y)�t/>����GE�3�9o�^>�#@�WHcA`�o��˴ܜ�����6/�O��Ϧ�C�4zB�J�788�\��5���H^����G1t�%%8= m�>�Xq�T����5�J��_�Y/&������&c�^L�ݖ=�|����=�I#j��з1V��2��u�n���x֭T�f�uV��b���� �[�y[�[��I�#I:̶������ pb=Ƒv���CXe{0"���F�ϵ/�b"ﱤ��nwh�����F"T��I�|>D_�}S��t������=����,)�_:�T�&I�\��@�d�UL8��n�Q�w�88]&�܃�{ެ2�Yp��o�Ї�R̶Bvz��06M%�Z�X]�hgZ��0r���:TS�k����J��. f@�i-��[�6'�����*��iD;6fwl#�W��u��4��#���v�� �]�-���RD�VQ��Iâ�I˻!���F��ݎ��k�4�q$��9b	�ט�v��u���:Y�mo��]�ņ�+{(��ƶ�iW���%��E	� <{Z� � _o�d��^�����J�+���0>�e�l�F���~F�8[G�����Jb0q��������҃[�振����^�Z�������,9����G���ۯ�s:���f܏�Ʒ���w�c�&�m�W���׾-�A8PA��w�>L5pf����-��&Q�Rl�TՅtz*�{�
E��=�
hYݭ>�J�Xn3�n �j����Ĥ݉�$i��F�7ͼjy�&/s	}L���� �6����Fix,"bN����ٻ١�G�ID����8��sR���(�� �!5�M>*�{�w�f�]�ő��i��Dٲ��ĉs��>�cݺ���9җ܇�[Q�������1�K#��z{f���C�e��f!~&�}������<�q�6�4f[��+}��~�K�A����H���F�$Վ����J�mt���{���vicw��g�j+�3,����m�;Y�@�=���Y�����!�ъ+e�Iս�Aw���7��%C�V��l��_�p%�C+�ׇ�{��bFB��J-?T���]��;��n�k�L��28|	�S���^����hQ�No{��������/�Ck�ڪ�����������V�DG5m&]��5���MW��=�P��mj�:E�_z�&����4�d`�}�[.{�]����лҁЮ!FT���$�R~86>0�bȜ�K7�_Ų�'�X��}GHIr�* qQd��X}�`IZeBZ��0��r�'���bmQe�6��!�_����<�Yj;��*[F�dD��Y�c���7�\M5U�Y�Z	F��k����h[b�~#�|_��D���4W��i�n5ޛxL�߀�,Z�����\Ф[�����:��_���s>����xJ�٤�B�2��#9��;�R 
)�z�|*=��*�O�'������M�PR�t��Y���==|mЫE��J3`CΫ��e0���>dY�~�f�ل[u��MH�Aܹs����Rp��a��6N��.@E)��K�<K�R,]Wԇ��'���]�c
�Ҍ�Ӟք;tuʯg��(a��^O��y6�J\{������	�v1n��g�9�	:�Ca�ǉ�oRP3+bN��k��	<�@6�eyN�ܶ�p�=�{�켺����$/��f��slF�s(-�%"{��&��pp/Q�Aͦ�\�ǟ$�a����r�lX���X�Tۧ�8��pm^�( 窼P�P�v��I��7��K���c�`O�%P/��f��z�(��&̮JF�i�Pqc��;��#��L�hĊ15�d�\-F��dLq�V�����b��\���Z�X�d�
��ߝV��,c7����ꥪЮ�_ 7^�1Rk\eX�9<���,��f�]�Y���e{DkU�?�;9$���u[�S�Ѿx?#���Rߡb]X��h�Q{}J���pMQ+�0�!V���M1e�xZ��F9��_����gu&��^ �e%��;=iTƷC��ߊD����u�]%5�S��/�,�My4��B���wS��|�$ (K}��3[��>�υ7�:�l[ Y ��p�'H�]��&)�ѥ�=��h��Oș�B��"����� Tw�uۏ�9k�=�T@��^�Շ%��ݍ��o�[�]�q�A|��jO���mvEZb�*�)���V�~y:9 :� ��"y��L����V��uZ=.)b+�m���Č�b%'a��,��,5k,��#�7�k�$�mB��JvJ��">�c��w��!+/�!�?~5�8*Җ�n ��B2�?"���C�즾Ղ�������Z�
f������̅��G�pdptd��@
Fn�
�BܜY�Z�5	;�u�����X�j�x^؀W�~�@de�>�bߋ�u2,��;J���(�Na�ғ
�Joږ>����͹w��� p�=��}f!�-�T�)p`�`�)t��� �}�E-��<��V�`&y���0A��5��V�s�B��j�ͺ ���������c�(ߊ�n��/r�e~�* �j^%�e�dQ/�!����[��t<G�B��kҲmP�YiH���L1M� $��}˾ѱ���7^o�@�N�(��Ը�b�X�^dYz���{���L׭�y�s*��#���鐎�i�Qgw������/�xyI�ũw�+?�|&9�.\���kA�ʡr�>�K�C�_�I>�49�#͟T�wDU�A��I^����Kz���MkF���h;�y�dE\�P"�X۷�>�o G�:Six���.\�5���u���:{+C�[{�~y0���WJ�u��эd�U�T����	�k���b'��)s���N�`�K�ۋ����0��xB�;V�
�\��1��[f��mrr�`�b��t��%y�6�u����V�(��+���02+bM�׬4�8��7�.a��U�$�$��~0D��=IP��K��1 .V�'i`hb�1=9�&!�.��k��7^��B�fT�<�����.��}쎐I�|Q"���78�3C}���_כ!�����,��w%8% ��{?�Y�$�cUL�1�\��$��:TQ������&�����5=iO0�C�K!9Wa�IXҽ 5k�Ȩ�<sy���tյ���	���T\��E|��=3����^;x+�ߵ�=-=�FJq@����{s0�/?�����$����ל4M+�~y�Ã�[>�9�,ޙ-Ќp��[@S��=qE�ˈ����ԗ-���1��D �0=��]`��t#�z搛�܍�TM!�G���,�fe���P4��GJ�u�O62zU
l�k��4�Y�i�C2u��jH�s#��qIb �5�i�4��7�i��Mh���.���s�T�px<�7�V�=�}������MQ��ȇm��d�S6�oR���fl�!Jݯ;�Lb�HP�3���m".�N��8E�D*��Yx�t6��T
��%�]+�����s�y�� ��l����#l��ؙ��;~a�oc*�2��p��Qs.�:Դ��j^�*w�I���ZV5����7s>I�����]�XS�`�I��DK�"����5�����D�Fa�-�-�����NY4����nG51�IE���Z�Jl��"��/9�6KL/3vJ�l����S�b�N)4~�6RL� �5����M f �D��R���܄ń5��Q�T�����3iG���P���۹.�ap��uT脽��a��sz����d��w�.�:���oA��)�B:�tɒ"$K��13"m�%	(�G+��2�2�E���R8�NE�(.-}�O�PG�O~V�5!��Tl1K�N��4q�"�{��9r4߬鑓h�&xn�,�?خ�p�3C�]|
.L\qtCO����J��n�N�;�'�Hu�ۛ���霨���X��ŏ�.�0���H����ocF-��	oc�d�e��p�.�$]�~�����Y^����-��XioW���G�����2�,?DdX��Q.�����Mc���6�$�&'��
����%�­?��=DY�٪.�6��*�U�d}l&tUf
`���C����UU Ibt�� ����}�C&n�=A�:� r1����&j�Y� Aߒw#d?;Mc'"��k���h���v3G	�S��q!��K ����m�է�8�֓K/0��3(���ʮ!p(�f-vD�u�X��l���:�^ ���z��vÆ�����e�Н��DFԢwm�1�aa�v�e�۝��&�c;�����7��!:�"�]��$U����c��a�{{���b��������Ք�q��Z��*�q���/��y9�9���$"��Df�6��P�Z�p��3�� D_��	���I�xq���ޤ S�����i��,6�=m�XF�b�����>���t�+[����s���/�NH��4���h�W�׃�)�Ԣ�����ۆ+�u����R�lQQ�ɩ���	��e"O�|��UH:��N����|������zj$����y �/C�t���Hd�]�Zpjо{#cc�?�$���5a�dB�%1T���cU=ũ�r͟wa�X �l�8�R�]'��"�z���V70)�_�$L��s��nS�%�ڎ���ڕ;�����48s��L�?�D�c��������~�RHär=x�9�g
�ꡫ49b�r@���"�c��=�u�YkW�hO���o?�r+ ��KHV��-c>G�>�8��5kÝ�LR���]��&~�Ȗ-��f���(`�Ә�=�v��:�b�;��L�j�@74�W��̣���x*��M-��w�n�|�ӌ��_�&�οg�y�B
���/��r�~�͞�x`�@��J�9�i�c�����l�c�\��l5��<��;/X��W^�a0�Y x�F���`�I݃�[�<�z�#��ѓ�ZLg��Xm�Tڲ��̦�r7�v��Ib�{�Ę	����눎0�T��#2�Q��BY1vVt�� �ty.H�ݾ���� �v+���Qc[�=2n)=S��5��!և���MFs{�P�%�j��-0N �:��a�⠶�rY>UM!Z�eC���
 z�/�{ġ����2138Ok�
����̊�����H���a��sU�n���r�&��Yݔ1��耤�Jw�x�:��}B��Qi����Od�)��O��=���U~2�)Y=�C.,܏��& m��6�<Z�o�2GZ"9Pؐ�P���ɉ���L�#R&U��C��u����<(�IAխM�ٴ�ݩ�T '����2;x�$��%K(\��-&|Az��6�c�s�l<V�\�;ǦA")�(�>9,�͞�%I)+m]@�-��Ѳ�6��2�Y�3�j����|�."qV��ۡ�x� ����1�>"\u��Dػ�c�>�
�N�<��T]S��{�TBJ���{��x��
�
-]Wq�y��O�W]j��K�b���Θ��h�B=/�����C��!>ˍ�r�hP�hՃ��0��D�*da��t���5���M^����D��Q;�Lf;��O7��>u~@y���Ϸ�e�T���e��/�=�79�l���nC7u��������U������/腱�k9���b��cr ���I�*9�`kV	j��O��x<�ʙJ���+��P�?D����������N�}����-Ԩj��8w��ؖ:o1��tS��m�'��XƇ����e����{�!3��C���UEOJ�g��A��Q�zT�,�x��H��t@���n�1����Xt�,}s_�z#,eZܣ��N���&�u���h�s�5�-S)�:��Kvt�Mx͂� K��I����g�˫�#J�ee`�E$���}щ�f۽ta&N�R볡9i���r�v[bh@��n�>k7� �U*S�&�-�un	���Ƞqm�"���8$����Q�I���1N��e�S�]�?F�4|�:z��x$�W4����%��^	�*:�?E,Q��Rg��1��h9�5���g��@��,l�����if}�v�J�Q��`φ�	#VpY��^����]�'�	`���"o���c\@�ק> ���t��W�{?�@�ʟ��D�ʽ�}Ac�=�$e<�s�/@��!-���*ϲ�4.
g�����gټ���n��Q9A��r���q��x�^k���`��������ڑ7gPz��n�ؽU�У|s� ����1c_�4�`#:j����r��+@:�U���=��h��fH��dxBF�Ͻ�9�o��S�W���+)�A�a"ԫ�m}�j7��<��-��	�EQ��w�fS�m�Z��r=֯F0��t7�mq���5.��N��,��d��6����h�ƀq4M�BGd��/��Y�-K�%y-�O� $�OR�j]y$[�V�7s������Q�0��S��v)z��g_f�L��S�����Y�����hu�)X����\�GeF�� ���]0J��9V�x��Y0�~S��W�V�l����EdR�/��!�_n�2�)J���i)���rD��◹E��p �n��wo�i�6��o��?����	i���+�n��
J���ą��&��b@DiƼь �_�ʆ���֔����8,橋y7`��#�G r��b|��|V�+��g���g�ڂ�μC6{�Z�q�1%�Cа/����(��9��z� +�F\-��C4P��?۱��{�,5`D2��t?���V��h7�0����]��/0*|γR���DƱx����(*A;"�*����N���y����h8IU�6nZM'ʄ�l��;��}���B�m����8��an����Q���$�Lr使O!�Z�5D6�qg�w�X�|�fQTѰi�uſ�-�R����H:]���n�A�M4;�(p��YD����9��q���v@� ���{Z?���I
�0�+橾f��H��T�������Q������4]殠���t\Q*O��'�NǪ�a���>V�澸�`SVگ�����/6>P�+fz�:^>��l0��Or�Pa������B��ՊJb��CfVm��j.�I'��.�5_Z=!���1�G�~�f�H�dw���	��&ߙ��{��g�U
"���Rۧ�N�wq�(<P�acaU{�>����[�j���������g�
���ϥ�x���7�_;Q���q!�K���̚��cJ'B19�R��p���)�w�[�$�b<$ik����a?�\������=@0hR�->I�UZNt�ʴ��
_t�i�kñm���ga�U|ӘcJ�[V+�B(�%rT������i������לVS�(����i��ޏE��z6�{X����A��F�C��0���+Έe��~�D���Oqgۣ3��8MCWU<�F���k�scf�����<Z�Ki�v��QB�n�˫���ϙ�'��_|$ 5�f���l��/�F�~�@�Q`pzsT���V�F�y��lfN�U���p�P$��S���[���2����U�p�Y��[����b�I�f����:گ=���+"UM����uo�J1�8����먺����L~�i.�GH��pi����6��-x���pPZ�$�z5��T�AL�p�%F#�����_8m���� ^يq��3}��Į?h��*>�hc�R���!1��Se)���)�'L�
�W-�t�C,NoeL�ZԸŅ�`���
A��Z�s�%�/,�G�¬�`�  Z`6��uJ
������ûh��s�C�DT:�sڿ'm7��n<H|G���T)���~E�Zq�mT���٧9��ʬ�Dx7�����x]&*��Ƕn��f��7c�"�8jR��w[m2���O(!�Uo�q'_�Y��� �)b��H�%�g)�m���q�4t��*�W�Gp�tMI�����<�5]$ؾ��b�y��w<�❿��q3z��x�ਸ਼�Y)��bԅ�-�3D�������3��3�L��]%�ѥ�Lw�mD��9��c׬ne- O�QRH� .�Q�?j-"�9V�^#vd���-W����Q�)�}�7��쎐��7A`,��X6�`O�/敺�4&�i[	�C�@=l�͠3d���B���6i7��'qD�t�*�}�+�u���'���J�7�ea�h0�7��r-�26�=bm;h��?d����<5���\P�=SZLk���y�"J��r�>oo��-�čc$�Ù�A�R�=�Xj�s�橇�A� ޱ����'����@w~^�􆎃:�B�	٬)�.��Y\$����>X�ʑ�&��b���Bp�2��*���S�_@$-�jb��f*U\
�B�ƍn"v�SqV��&ݙ"�?�� ��;�$�.�u�P�)�Se�^'�H�Di:���zݥ6)��wj�[��Kj��r�Y�dw�f�ZR6&������\�{�l_ۙSdW:����%���)8n~�ق�Ηj�k����[e��:*c2k!�שw"�p@�Qz��)'r<�-%|�� �M�i�&,�~��c�e��(dvY��t@��/I���*+a���9y"�O��W�M�f%�M��]��6�`�Nm6̺��
�����{+�o�Z	,[G>��"�"��E[����P�����U�\v���s%�o
�(�bZӃ�R�8��t6��6�~ �!��=>_^F��:)T���c�.^��"���#��Vy�~���ѥލ�����'�D
 Z��~�fŌ%�M2�2*�Ys��u�[cao|͇�p�������syKF='��,6Z�dZ����i�#kI̎���h����8Ci�#�|��ziͱ_��C��'�V�O��^A'L���5�H&�]ޜU���W��&�Y���>�ƙ�h+��0�U#:���7�7��4��}qd��<�ڧ�nE#ψf-d��}������ČߙV���.��ܺΏC�_������0���I�"��o�p�hI��0�1�����*	�\C���V���E,�mТ��ˇ�%�g*�ZۍX
EJ���AT��W{��*�_�ɤO��Y`?tz\zӳ p���ҫA��+͗��8��l�����CK�s�pl�e9<C ���Z%� �١���KF6�l��
^�f5f�����〷C�Q��~��s��/wQuCČ���s������ÈK�(rMޥt{˗�^Ϗ���k {E�Ƹ�$��<-���(w�I���7����[w�v�@t�ݪ����WX��Q���X蠫�J>�Q���?���Waiy�k8��G8�n�D�ifiI�yy�G3GHx�?�G��.W��0a�N�)Z~B�*y�H�^�w�쿷+~Q���x���:%��W���4�ƒ��
5�����Q��=��,2���Ka���qW7��{�ں��a�ڳ�����ₜ���ǲJ����hW�д�"��n��]�����.��b��e�rP��6���i=x^t1���Żu��P��\a��0�1;��/+��>5���뵺���U��Όp��-*_E�]���������b��`B��o���u�Ո{�>V?er}\msI2�tۘ���@�� ~G_>G{�p���Ŷ��V0I%�5g_ß=�uV��9C�QR�~�W4[�^�Rp��8��̾�~m�߮��e�m�\vZaDF���z��B�B��wѫ�JL6+\z�c�'���le�|�*�8��c��������'ʾ��fv�c�#>�1�&*�̟�"�Ś��'�������ON*�Ai����;�P������a?^~s��[א��ѝe��m��/����_�6�@Q|ժ����K�	�n����Y=��R�ۍ�7�~^~Dc%�>c&��ic��?}�_��6��(�R��_�W�]���ȕ��� &�+.�$�F����JXʎ��"|bԴ�{�3�R���u�(�+�9+�땕� �UGI4?O]�,��%�w����h��U����6����g��:{�(�M4��z�EZ0ma~C�i���a"]]P��P=�^��M�5"/d'�M����$����\�S�b���;�X��X!��TX���; /��5�#��on�h��E�����C7�ӵ
�h�bk���=s�#�{�Zt��҇�7��to�s Ot�s��'u��.��?$�.���5i���H�P�9�}tX�-�&�O�6���ɰ�/׬v�iX���e��?��]~�����iH-.́l�]*P�[�Gmނ6g�+b��E�����Լ�f�27Fg�H4���A	��T��g�>��f�����!�i �M�1z�	� .D_��U*S5�X*�lǞ�F��p�%t��6=���'cj�l�n*�ýs��N�l$k}2@_�Ki�3n�$���6�9{W�Ff������.H�Ђ��MO�X�J�{k���8Z][�i�/�{	�	��f�yTI�
�3`��ݼ����~s�h����
�$��z�
{�X�6/��]���
��%��R�2:�HP�Qn4t+��_��@*��Fnr�u�^������ݲ�Ҹ{MS]�-ЖF���+�y'�&dk@��91��-��#���o<AA:�
��M�wߓ��A!����D��HY��e�� !�&���� f���Uў�.F��2��m�8p3EIP&���������r{�5��Y���7	��2�s�j�0t�2a]�f�r)������gS>Φ���8��B��@�^{pB�"3����$��9�ڔ_F�qvSe�(R���<�ԇZ�HL�3����2�����MV��f��j������b��$�P��y����V�q���L<�5��A�0	܏e
a��F�t�������2d���=`L_$ ��
Vkb�v�~�F^�Y�%r.�^Z"��4$�|�nA"Zc1�MM�����#�K%"X�'�K��!r1+�.f@��%��������D}[��fD�ջ=�5��� �����$bE�f��장�H����)}a���7� |,����u#����<�%S���UiꦙW��lo݆g��΋�׮��3��-K\�D��-F�k�n鮛���Zvj�I[t�{�a�D�o^��FLL���7P�V��]�����гn��{C� �Bd��)��Qp�D��i�g�٫��g��P���nF���ܦe�Z�gPa��	~�Ï��b����|��*V@wg� �P?�iIo�����G}�{v��|����B������-O�'��HP�	�4�@�;7���?Ϟ5�B�h�>YJ�q6o"|�ұ�	8�o�&'��S54��F���T��2�V��������Oo>6��Aΰ� ;��[� ~ߓ���
?��x���pT -3r�����e�E���61���v_��lԴ�L7;����\�K���D���y/�M�<i����z[=�޹�6u8,Z2	ئ���!Gn�d+���<���ccr5fV7j���e\񡰁���w��Æ��>��Q�������+uye��h���ie��.�	۞����P�_�!��AiBS��ћ�/ϡ�E)/�kFiW"���`�6������%�:�nν	�	fG�Kרĭ�ڿ���b�<�Q	�CK���f=h���w�J��-|9����ZN�����v�A �f�/}:5}���Ti��Dc�ҟ���E��~���`06sVS/F����SH�j�6����a�#��-�F�^K���L�D�ڥ\PE�1�~"M[�2f���eF��R��4U���i7R�o /�"��c}<�c���b)Z������)|v�e ��GJ"�"-&3F���c��A
��т���v���T��k@.\˦��̕��8�b.U�ءҤo�����[��T�D輢Q�i��f`A"΁�ھdёj[̐�r_p�
*&#�|��烉��v/�e"t��L�vκ�D�@u&�ؾ�_?���z���¢����[L���h�Y�U��G��L�"̷戶(�Ҭ�Z��������n0a��ݪ�u~������܍��M,��p�y�ٚWo�%Őf�yj��M]ɠ��wX��&���Ũ�7?!���bc��������ݎ��L<XK���(ί*�c�X�{)�m��=��3",]c)��l>�Ë�6�������J!��m�)	����L��"d>*��$��%@�-]���L�޼�[]�컨��z��#)|��ٙ8vnBbo��@�*Q� ��	q���5�P6VR|#b�̪r�M��h)�J'��6$���-Q��:�4�O��_�g�YY�#��0�=�sY0ִi
�L&�����(�ͪɁ���@<��J'W0Ӟ�#z��q+��/��	M�:_)�����,6���$Xq<E��z_n���t~ĉ�n��p9߉$����QL�Q�,5�tb�O.��&�$���R_S�ް���K�Ŧǉ72/k#j�<�t5~�����I�r��[Q�+�v[2�VB$���Mv��c����O;��mcFR��3@�hz?Q8DLb���>���j\����~L��-�-���+0�K3��:]�~u�?�N��Ԇ�#������s�ILܰ���
[�i���Cg���x'Br��v��5��͈���PQ���]�?����m��Z�`#RaW�CS��@]N��*��Kĕ|P�Ya2 ��Q�|ᥡ]�1�=X'���_7�_��ruX;K!����R{%�������O:ޠ"�"�⌤U��,����w�� J�H$u�ܧ�3	��΢���d���|}�6�D**^��8�9�cu6�;�w�ǜs�I���3=��BN���hO��}3�<�t]9�k��Q��{#��jb�=�F�o�?�w�������<�D��&a+輧�M��".����Q}��<�A�`��o��)�l���������iO7|��@�O�m<�IR�|��u�	�c%��
�-������C�����=���[@�����Oƈc����rl��L+�@������Y���5���*R1�����%������� �����kM�8g�G[���9��xa� �L����q6���;����nf{�[r���>L��Y�D:{AZ��Y����k���T�B��ft9��6_�J׊���� '�jU�]xtu�Ŭ$F~�ВbrD(.ú����R����zQ���E��J���5�!��AR�%	vj��ƨx�C:��afNS�������T
rqC��`���N6��*Op������ġ���A�E::q��v�x~ ��\\3��8O�����M��7Mr�GGr~2~�Lq>^����Iݜ�0���?q:���VࡴO�KMVߺU�~d4�:�^�E�m!�(����JM�����u_�1 � ,bh�Yh�������]Ճ8c�\<ŀ�7G��.>�A�XW�\b�..��a����o�,�sw0-"��"E!J�����Zy�+F�y���v����x�7��`�� 0Hܱ�#��!Q�q��8O�wJ�i�l��Y�;��?f @(bx�bJE��r���;Z���05��c�Ce���q9%�B�.
��,�>Z��F��n���-��}`y9�1 .ˣ=�R���JN��qD�V�S�ğ[ƃɕ]����YW�#d��a@�}��e�<���:��/�Xq����a�L��K
ɱ�6��4��equ�%p�WZ�d����F���HU	Χ�`۷P����-��OU)/��M�_��Ka�4�����*��s�f0�V*E��*�x��6?���|2�6O9�ZQ���۔hJɠ8�ӓegc!�j�In���ܼ<�X-����T.�_�ͱ|�l%KJn����m\����Z\�j��GR��b��<����oo�RDn/䎉<�1��*m�Q;bƭ]:�T3�g�qWJ���De4 ��ޫO�TJ�\S��0�=k*8cy+�keoB����6��#����s�B���������X���Bc�\KJ��8^�=�R+�S�.$(\C�`��K���%D������w�:�!17D
�)#Ŝ�r�fSK��Y �I~o\��k�ב�����>'�o�(��Ѓ%hb�:vo�[P�n�\4~+t��72o�wtB�T� @^B���#��	�t��]�}�:���a ���G���4tov�rLOr�X$���f�:��Ȃ̵�~�Grdު�]����$<Qn��ɟ*q��ȕ�6{ȯ��D,�݁_���È���BJ�h��D�
������M����2�f�����r�h��|�Ɗ�ɜ���V�����G��p��޻1�S9zHԃ]�6�B�4ٲ�ӎD̛�M��Ì��ib�]�O���^/���s�8�/H%�-�֦��
�6�T����z�R&������Jڄ�����Xr��Q��h�i�vzI����˸�W<��rX�?��sf2I�c5cy�i����q�#=���Y�鈻�>�G����{�A@ፐ�k�F"ԇem���`�|RQŊ," �$	\Fuj��ϝx5����V�K�	�G��W~�ȸ�.�1���9�w�-�
1�������cj�\h!�p��T{K�����6�I��e��E��@���?�65���g�»)d w!�����ŁS�%7�#�g?��q���G� c@[�T�%k�մ�nʍ�^U\�h��j������u��E]�.:vWsX����]A�p�S���n&�gW�d��4������fR�r���>����R["ƕ�* ������)���|�����#�������G-wߤ&
�Շ�$��D���]��<B�����v�m�'c�%�N��Ԗ�ϥ��썔8��f]bח(Z �@&��ٟ92�V0�j����ۚD'���/�븒6�Қ�KIf��NR|T4S�a_G�6/���Y�%k\����z��ώ�,Fɯ���!x��5'5M�':1w}i��nG �-c���ȟ·7��<.�Bo���^	1���~}b\�F�C��Ʉ�.*�K沽����SS���bZ?�u����5��P�&p�:�����Y%���6 ��w��m��Ɉ��;7_6ΰ��>��Ш�Q��չ��WHE&:���=ԋ�l��2�� BhM�!�6�H�efL ʎ������CÀ�e2��l U�hV��Wy�4��;{��]#������{=���W����BChI�\y�J�ް!�;��9x���I�㓚�6u��S��U>������ �׼�в���̳��M
l�%D��y��*��_}�!h����#4���1]su���~�1Ryj���I����7-�� ���	�L��C�z3b����d,�<��Ɉ�0\7�7nY~�է���� ����8�=�`�� w� ��ϊ���c�����R=�(M2	�ę�&���v���b.�?��6�pcav�AU(b��6N�h��O�~�mw��R�0���`�Gj�Q��Ǆ'� z0:Qj�
�՘��&�D-Х��('�7ߪ��/�_,�6� ��I����xm�u����ae���h+5����P��ǯl�8s)��q'�T%#{�T�����g�%d�����'�}�2���iw�j>Z�'H��v����j��콞!ڊz�tZ�|#$�o#q��iG�'�Z�$HR�Q&�fsu��j?t�֐+H�-[x�m�Z
A<|��f��s��ԯ`AZS�;yv��rڑ�z����E���'�l@���h�z�J��a��<�Z$�:�<ß@W����4;2�3�?)-��� �է���莒��Z��@p ����&Қ�1��F)Tj
�-��>����m��?��Wj�͂��o
�_;�p)g�(]�&��xݒ�n��ksa#�Y3z�f9Vԧ�<b�@�*\��c���ݭ�}E`�k��\��k!�J�#�+ �H9�l�g-�
Y�1�x�f r��$�{13)���T6�D�tr�t3��于����J$�w#˽��2%OYf/�}�V�9�zG�h�ɶ�LfDn�/�I��|q�hS�,E*a�SL�=*T�l`}��n7��K(5�`FL�� ���B5Gɠ�~,��������{�I=��ƠS^�J�6ʫ��
��3���g�	Ǌ�QS�R���2S%��zN����IW���E��#�z��g�>�G���r�?)`BS>�
Ҍ���<��5j��E��>qbi��ï%y�x����^tU�1�����:�=�>$�:_�<ue�ƿat���`
�b?!^L����W���K,tO�<�}LD�yȔ2'�7���	hJ�������>�/&���(�rƏeʧ����w�-tTPL�e����hԯ4I�yAJ�>fK;=)��a@��|�j�v7 H`�T��JB'Р��U�3��1����F��3=��>WilnN�k�j�<�Nkp��l���Z�0t�i��!Mn����T���*{��ҳ �i!�X�G����&�����~�R �\�ZMW;�<���A)�5l��=a�t]�;,*me>w��z螸�L�{5�U��R4(8C�e��w.�@�dQ���Ġ2��΃K�ǆ�a�I����f�:����%�� �!/;	��]�
� �; 4K���EjGs1_�����g9��B�hrTN,��q�-(C���=��ڎŻ�*EX�y�V���W�N8�����>lJ *��Z��"�ۗ2��Tঋ��&�S�ēd|
�C�=�E�3�ٖ�L#��[�K09>��Q���,�����'\Ly�W��j��j{p�<#Q�LX����-�VCl1�HΝ��)�Ƕ�m���\�0�uQj,��dh�o�?En��	��Y6�AO���H�R0�i�a���bX�oh�!��kP��E�H9%,�8J2.����of�y -�|ff��:�Nw�(�7!_q4�z[�)�Q�	MH��0f���# �`�z�Q�3�֎,9����7�x��E��.�	����,��kM�>E=۫����?���p�x��I��<�ޮ�P�T�TE���k�N_�+������.����S
$��|�Apw�s��q~v�s��п�S1�W0�i]�V����D�s��a�����2T_��Z�L��ؾǋ���(?�E�p}�%�w�uo�a�8ӿR��X*՗0�8E�e���/ſ��C��ν*�#׍��B{�;�qM�{���k,�Ow�*H�k�z��`�٧�s�^�BWB!M�|�YU��nՈ������v"��K��8>�=W��:����6�#�!(i�丼�
��o5�B�<R���0�O82Z�äV�^N�ӆ����w�-�� ���w2!W�B�a�����.� ���;�P&�ϓ��s�V\՞�C��[/�2+�샡�ZF��O*z�3VC��L���`����3��!C��$��U�8	����ͽ�&�L>?�'EOP�|�S�5Lҿ�{	n/Pfn�?PM�\�o����7D���7�ۈ:�L�<�+&B�ҨԞ�Nٍ_��n-�����B���C�L�f{\����kc! �s��ڒN�?��n'0E�!�HsL/�[����X�!�<�V�x�+Q���o��b�la!C��n�0ݏg�O��7߿|���0���E��t����Z��R��(t�6��{L�s�]MJ�����{�/�W)�Nk��'��X�J=�
���0�Ń���$:H�@�hg����*�KU;�N��������FM��c�ʉ_�D�Q�=�an�7��3![p��jC5i��&bPl��(�����E��ͣ�z�����t�����8H$H������4�Y}Z��g��u:ԡć"*"�0{�f� �����B֙�@����Z1e@��a�0ߞSŃ��j��Z��5?��:��	�vl��A@7o��d[��bJL�x@�o�8� S�*���s�.�޳tX��4M0����|N��H]=���n�,�WS�ߗA	�ݱ���T�����ΰ���[vE�Ƒ���q���K�i�X{��I�Uɨ����`�{�5�aK`�.�Oa��L�_sE�B�_k� ;�t�]>[Ȇ܀���x�{8ըbv����H\.8VP���eLg3��*���2VY�|���8y���q�E=P#y��l�-!7܋0p���'�%[(M]�=���d�!�S�r�Ph}��EF����D�<;)!�绎>���mY�b��C�P���֡���,�3j��%l]���^5L�]y�A�[[N<$g�O5/��>А�MV�p=@�5F%�(\�[i�����K"��\��ވ����k>'���N^E��g�������E���Uv	�B����hf��uO�`K�X����(�V��K�Y���Z]5Bg8RA�ޞ+��Ļ��2"�XA�_o�
F�:��fZv�-EO`�w�mvl~n�>/�5_r�0�g'���Ab7�r[M��;�C/�80���n)������Vu7����Yl����"eȥ���2���AXRL��U:�;��+[;�ف����$���+u�Ԟ�s�":e������Zn��f�Uo���Hr�[8Y��ɵh�!&�Mwx=C���^�l�U�������j������s��n�����[�'�&���,�q��Jȫ�wĀ�]�Tg��j�Z����f�4~W�^�_J�J	TB�ǜ�(�:�r���,�+0��%�^�R|�$��~�*�B����9P�Sw�AT~]����̬�:7���e���x�x�Gn�)�bћ1��"pf��4�&wS �Sb.(���$Z�b3�M�q�/�e�8{t��E"]籴؈A�gF��x�l���8�9�&���I���U�&�_ք">e���^���e�_IV k��l����
����Y�F��x�/�A���n��o�3���[��	���^�����%�wǛŗ���3\���k7 &D��POC딓.(;��~�mv�Eu�&�0��J�� �8!�r�LP�C���Ox	��T�@��t轸��vR�����"�UXr+L{x�M�z�Ybj}��1P�]rЦ>8�ɜ�S��ߌ�z��I��z��v���!B'�R��󔔌�a����(�LV�Ȕ�N`�A��5""�9����9�(IP�c��qz|�Mu)�6�����@JG:q�r�@wY%b��h�ܩS�L�m,�S�5R;!��8�Y��=Ƒ>���ʮ/ .�|0(?q��-�δ�&:�ܓ��p*��iA���,�z55���1�~
�b#�!{|�Y~<|������vȧ>7���jd���ad�]�+�&���GSi����Ц>��Z�\����pl��,K��;��7V�j��J��+(vŃ>�"hx�EW�bʙ��2���W#�ֱ덒�51!��V�[nfڙ���P>2k�Ml[�PA���c��Ϟ R�א3-�~����^�߃踌����q�R�	�ws9P�2O��w�z��?�B`3v��w-}�,�{aN7���<�T�y�H�O�k)�r���[�
�T����A��G~�F�2���£f�sƓ�d���|���B������,�)JTp"�A]�ci��ڨ�J�H�Em���Qr��?[0:�Ͼ��\��N��fwn+]a�!���L�����8bh��Ś�h���_��WN71%~���8K�?F���R�ZyOTt��8^	d\e˰�QƬظ
���[>�Z#Wf���\�C�T�FP���>j<u!Z9[�vy���	�|��.���@V���� p�d�� ��l������Pi�-o�)K�F,�|�XT�uė��M0mb<�M���>X=?�I���i��b*����3qua��j�;=�}��u�:�/�i�A�/����� yo��n7�'#ZG�s"꼢�WG�+����� ����T�����S�o,,h���n���q�Λ	
<�!X�'�w
�bp�7��.O���.6�XM$�-�f݆g�(���� ���/�l�p���j@�Y[W�NZ��� �y�E��6|�X�>ᙔ���C5���nG4ba\:B �&����z�"������yL�ѿX���Ty@.B��(����!�^;�[�분��K�\�?/H���k����ڰs���|u� :��Z(���E����Zi�A�:��Bf�ؙ���k��?��_�Al{)P��F�u#�W��mi`�]���3xX�`����E�y^��
&�k��y=�gǗϐ�~9�)���#���D���J.ͦ��{��}~�����(�u������!��>�P���gR�u}�<WN�4cVq��uJ�B���KY�e��'�=�	��(�$� ��'����б��~������րP�O�Ͳ����n�D�B���S�N�����$���m~U��;��Z���N�>� S�..X��;���DP�%�ͨ�ȼo�9H�*��4�K	�����-F��}� oQ�'@���i��Y��0�j�]!>T0��7��"����$4�Ke��������A�<�d������`�v�lӪr�ߕ��R�d�K����"���8+ï��O���v���Ši�BC�~�3 K�+�3YGG{]�>b�?�O3J��*tO�����%��{ 7,k��yWۤ��S�ھH����e\����)���� ��!����Yp/�m�~O�h��L2Q;
��n�S`��UpL�4!}h?y�Ɨ]ؙ�N�P�KH�3\B�.\��|�����?���2�
I��v�]����p����>��yS�V�Y�������n���ܬ�L�����xm@�^�P������5pS�^�잀a-g�շ��3p��b�_�O*��& ��o�4H��I�qհ���� ��[lJқ�����Ӕ��y�>_��lڥ�xy�c/�GE���vM�!N_���|𸧱�M����*�^������Yn f�a �����"F ���&��Ѕ!����0��%�q���1,�/f�m��;�]?{*Y�Q�P���(�
����=�*y"�M]�l��^��
ZlB�ҟ�^��.J�>ز qkD�P�M_�,l�,��1'�(Q�U/}%��n�I>X�1��sr��թ�U�N��¯E��"���h�]��q��Q��y|����5�rCc�n^���� 5���P������)������V�&��!��D��FK�B^��<&�S�H^zX��y�G/t@��~x���?��dZ.��c.7N�p� ���FժA޼pv�ߖ��V��U�Cru���������	��dkV��YϏ�%�v<�Ե�hD�s!������b�[-%Pb�$5���@]pFI5���E�m���G��g�SJ-�`�A	��iF��.DM{i/JV�9d��?��w�;#G�~t��?u���A��r��zZWH��]
Tu�!�J6��!К���݊�ꀆ���쓖��˟��Y���>J�.�me.^�7x��(�k�BWޣ��(I�Y�!�hm
��\@THYdxO5�7�Ä������0f�W�>�\�� W�nx���ۗi��(�쉫�Iw
����oh$!�nT�yQ��ӆ@���j�9�� I���{΅h3���}=�6�,?��X�f�Ok9/�n��ɬ?�ot�U&TU�xxi
��ƥ;��An�fp�_+OEpH=vC��t7����3��Ƅ������ }�L���<�����!k���/ٕ�$����ڄ5�bOu�Ƭ\���������o���z��Y?�	���!:Z ��n1P�-'���rk�i�~gX$>�'�P�Y���c>�ƣ�*ٺ�j|Rz�딭I�ʈ{�p�md\`���^��Ƨ㙄��~����'�6���V���v)�(v� ?�R	���{��&H��*{�9�[���8�W�0�5H�蓠;��?�f��Jrެ��������KŽBePC�P��9":�/8Z[%8�<�UtR��'b��4�7�ٍk󌬒��t��<3����(űP��N�N������~���EVL�c�&���^ ��`�x���I�����i�p��n
��ǋsJ�h����ڜ�U��V�����uT��x��/�$vgz�ɮS�Ѧ��cǷ���(�G�z���n}.W}����4] *D���TD�� ���L���~��D���\�l\53�]�5��������l4�H'��LN�햢:��x''ՅҀ�	�VY����-��P�?��� 0���vۂ2��l���l)e���(���Ǔ�D��k���aF���I{�T̰~�2���K ק����.lR�V;v�T�[�h��(\s)�xb}e�4=�Ue�?���ܬ��=����.��t��M�V���:B^p-~+�,2+? �4^��]!�ً����4�#'E�6��6p���-0��DX���������{��VN�?����OH��KǪ�"_Wn *洑0��ܭ���[���j��QGڇ���[z�IӋ��#R�9�q%�%��paft�]_�NT��jNa�\\=��-!�I!�AC�fRG�&�AZ����0a����,s�!W�e�G�`خ=�'�;Y���k��sΖ�Ø�,���˨ ���� H
�HL�ic��7���e(����!\�� ��i�xc��}�/P���a$?���MT}��"���8�b�/<~�9qi�Q��S�$&}�@�g4�@�3w�^8���]�-+wc�pY��[�J�H'f��U��Sē�oJ�p�*U�gʲKX-5Z�B��%⼻v�u�Z���̩�ҘV�K��)��"��_*�Q �z�D�Ϯ-��18.���tF��n��4t<CȖa����O�{�BG,�1�-r�C�m��j%�G���6��̉f�ƫGs�F�_���(��R}�ܘf�f��	0�Z�2��Z�l��Ix�0�W��-B������yY %��{
~����cdwnXe�r����Q�Tʜ�ng� ���eE|�Y\wwi��Wn���@��$r1�[��	S��1z}��ݟfcck����`�n���N+2�rA[x�5^"fF��Z�F���礁^цd�� ���M^M�R�#���w��x�H0���"V�q\��[9V)��=�B[�������,���y�s[�wqK������7���Ō���:��	�Źj'�Z�m�D�����Hɬr��-�".�E�Ã ;����G�emh#MK� ��d�zIQ�<�(m��љY���V��� �'nxd��ߣҦ�5�v����p#t'z�y�8�B#�6��8�Y���i�w���Z�Xx���o ��u�[X%̉i�9_����ϸ��Z��l����3�33TƊ2��"[g��(��3�3̽�a�:�e��~M�Z&��A@��q'��ּ���i��6:�8�N;�1QI1�%�_)���?��fϺ9W��n�q��9?ȏt�i����Rf���C��aP���£�"�U�$��ʻ�K��p���ȧ�2.Fm��M/�b�q�:�=��L��8�h���P�͘����D'���U�X���&CC�T���Aa<E��Fe��1�R\�m��yC��ލ�a�.�i�x����]�>��Au�E⽛��,.'P�+���:=�ѕ�m�8����E�Nᱮ��VQy*_g�P����G1�1(T-0dSRO�Yfn�\�C����W���A�O�&����2/�TW"5Xxq��KO��\@|v$�4���\"���������x���,��ԡ��ct���8�M�H��jC��d��B�+>�俀7��"|08&�%E��4�4�myņ��ǟD{ėi�����˃Ϣl��J��!7���ٷ��>8ɔ���/`i��:B8G�o��L=��<�"�vj�G��8�V_17�m=�Ͼ��(�j���T��Xg�iʳ�IK��T܊��3��N�$���K.��a�X��Z�����H|�T].���l���X�\�yz��U�����3�O,�?�w�Io&�N�7�*Nw��9��b�P��Lڡ��h~��0��v&{�q���%��J��<õ���Q�]jls���d"ɩ�����4N���A���eS#@�e���h��0kU�-�z~��E���ai��MObu���� �Һ������`n��q�՗�k
X��O!�TA�3M$���jdM���@G0�_g�lw���S��MO�d�UT�ăf̙��xL��y&,ީ�šSa*���8��؝�:�?EL2�4�X@x<�љn�}�5�2t&��=�q-K�i�m���Q�k�^��\�k�3�![�.�{����}��1s�W���9y��+�q��R��j���۠�[���oa�w۝yH�V#��ސ�������)��r_UГU)�9����$#��H<Ѡ��HM��3Uw��_-�EK�=����W_��d9h�6�j���F���^�v�V�N�m��Y��R7�:�UkI98M�ioC#K޴l��M�4M#���gs6J	�)�%����jwBx�@�SM��F�<�qɄ�F�OPzv����e��
v2�-�;�!���:&��"����s���$��/=�ݢ���4#Lࢸ�v{d�I\��7��ׄ���Ώ������wLLac�jlƻ�e8[-7����Y�h�e�ql�q���j��׭ը�]Z �L�/t���z���'3v�}�_��y(z���\_��G�@�'�9��uv�Y�â=tj�dƗ��o۹�NЮ����A�u���g`�Jn�yH���@;<�&�e+r.�¦%�+�V���.�B��\�D �>��oԆ���U�.22����1����G �9�.�_Q��K�bd4q8l6�n.7��y�_P�*�JM"�>ɸ�sJ[Ql���a�Tћ48�z�P�gmq�sY;�EZ�)K6��Cڻ?�a�	�ں���f�wR�ZJTm@��|~Ǩ~��7��O�$2��I{�����h��ΔG��@�X|ߓ�ϗ�`�-��+�8u-9����}�Pqs&��*�*U�:wP���݇��0��<PE�,M.�����Su���6Y�j9�j�O�����+�^�{qodTęy� "��-�s�ﶵ�@b�SI�m� p5|v�r��(��mծl�\�)�c����W[�
?�6,8=:u��Չ'�i;���ә���{��c�IL~�8�Ŵ �|o�(��P_M%¥c�W�'��ou��^�Gl���"+������_���E6�SҐ7N�vY|?2k�8��{�@h� �����x#��ƈ��1=�O����%i�$SF�)�U�
�b}H*U�����y�� }(�nG}�k۫I9�w���]�,9�2��u8��O�3���]�%J8�����6#�3U���AygW��8�}�1�+-���9J�BvVQ΀�0Y���Cvwͧ��ٞ=����+���
�j�T�AW�P�U�kb�qt]�c3�T̩L5�d��d7vK��W�����_�̘;�Oj�������Ō�|�HW�A�(���+t��PYD!�$�#���r�6��Me�PX���f�����B`��+�LT�0�&FgA��m�9/�a�BXKܔX*$e�z@}&�׽4���&Y���ufl=I.X��!�7�"��g��ҡ��|-�ڀ0��0X=�|�r6��u�h���B��×Y!���ʩmW[_�$�DwW*���0a�<��SLs�+�ą�b�e�[�ofS��2Z��c��؝��$�&���6��/�7�B�R��&����y�ΌW���A�,�@�s���3�ѫ���}��L�/w˜XV'�w�$���S �3�&Wښ��Q���m��Q��<셺i��ˆƜ��Jw�C�E\h���h��]�k�4���Z����`F�*)A��je� Έr�tý$s� �����	����!;`4��y�`�����~[WIr�\��ܞ�A��N,�W��Kf���-��� %Rwq5�S�S�����g��@���dcE�ʪogy1���~N�dOl�A^[s�f	Y�	E�o���>>
D��*��l$ �~�z�B$��k�Y^?��,�V��#wԘ�Uq�ۙ$�y�z�{i2=�f(Qg�(΅��8��%���.BX)S���`��c��ԣ������J5�t^�t�Dړ�Q��(]�|����vY��k�qy�sJ$Z���p:tH������i�P���f�cp���X4�F���5 ��)R��o~��`���ϛA� �����<���P�����W E��UB(���R*i�������[�����u>&-f��{�
�U*���3\��~:7ܡ�����	Qk� ��� x����/�]}*�W\�W����(�Kb$��?	�RD�?���
�T�K�-t�/�Qt|q�c�aR��xe�
�at��D"����_HuWh���6�{b7i�	�_~�N!��h�(B����>#�'ޣ:���Uuܘϝ�m�>�+���bR�b���ǵ���2'�,�����w�����l�j�cM��f�?#�`C��
�[���^�	��#�ߓ��<��2��̃Q��,暓\�b��U9��Cv ��;�gh�cJ��P�i��xaHI� I�j�� �^hT𝟔1儠�V�/�Ͱ���`��5cCq݃���]t�"�2�b���}�{o8�YF}�:1o�����"�1�o	9!K6\����5q�K���N�e���rc�{�^#Ʉ)v���Rl)�w%��|وﯔ�Z��5m���~�w&oӒ�g$���\S� h�K�ך�x@Z%��Ӣc��ÅH[��s<ZmC��kT8a�� X�j\�h���ot���&��y� �H�8��l����,*L��J�vP�Xൽ
w��R�����:d�*�|�#0��Ae��D�od���w4h�/�r�/P�Kzd����Xw�MQ/��}4ȝ�����W?M��`���V0���Qʼ�O�=c�uW������6EƹO�Ip5~ �u�ɪ\�)���jA1��hB�@�I^�H�k�[�5���2UW[��Q��U�ġ�d�p	��U_=��N&%HBw��~��d�_rZ���LW�<�����ޥX��%�����&�⢻�C�vRs���0*�U3L���f��I[@������y~dE0�S')W��'L��iN).
���^+\�l�g����z��K����Xq}TVԮ���9uo������"U�@�V����X�`�4�8&)gH�ZfC�"B�(/8P��T{q#��u	���,�A3��3q%��/�4+�c�"�B$4t.I:���k��:Z�R'�dy�E̛��!G=	�8%��פ˂�y���w*��?u�����Yz���he�<dK��C_x�oʃ��2�󇏋���4 �`e��L�W'S�2.L���#n?��a�g�R��y���X���y�܋bm��K��{;xs���t۶�
B9���!i>���`��v>k���)��Wم�w��;�r��t/=.�ʡ�£J{�_�(S�:���j`�[������*�H�#O����_Q1p����x�k���HC? �r���v���(��X��mb��#�� q�A�5����̫�$z��b۷-������!����Q1��~M|j��aq��C�!o+`�v�� ����nb�� krG�'Y�5��SR��t�0,�����*:$Q�T-��\T^]Z ��W��|�D2�����?DOQD5�/�h�	�M�+K���k�0��N����)�a!M�!�ǧq5�,��'۰&�##J�;�6Oe����#Z�jʼf�!�ES��V��]#z��	�S�eJn��؞��x!�U��2^�X�?�)>��N�ܹ�s���Ƴu	�>���%	��I�a"��5m�r�|�9]]\c��
VT����S�|�'�hʑ���?�9��s]�a[̺y&̂� �"6�X��a��^�����53HSW��-�] ���R�_�>R/=V�o,���b>�깫3�1���:\_P'��\��
H��⩱�$���H�UK�Ё��]u��*�ƹ�i��ī׏mϵ�ȣ�Ece@v�����7"C�o����?�k^!@#7�ҋ�
K�,D�����`�1�[���qҗql;N2%L����7aH~x׀Q�0=�(�!>���� \�j���;�HLLs����Qw�-E�A~�;b<@���-�����5��Ƚp>�uw}�DM@���xK"�%ۧw�#��}��1�G-��J�hw�q
C�܊Z�����ߓ�O�z'�ʓ����*x9�hi���T��E �/�}<�;+p$>�-�/��S��@��%�#�$����By�e�Kra5�u��xr�=���	a{Y�cT����AJb�B���!�򓷰K+�Hf��!Hr3�K!�(�X�}-�x| j`����/c'I��#ʇ��b�~+K��&�����-� �j6����݌�g�A7M܏��'I�4�W[���X|b�Gz�UL;l��.q%���D�!�S\��:��O
���WtܠT:2zg���;�%#��1��p2�@�AK�lr yL����YN+w����)��b$�������j��<Q��na6s�s�`Y��P�&�d6��ۜᑏ>k��=��J{1m�2��FԔ
����\�l�rp��
a �{Kx ?�'!�Uj�O�ȡ`,+���7x[Q�)
P0΀%'!-js���O���@cE2�5	/�-�ċLm/ 4��FF���eB���0}�~���:�.v&�F`Ar��ɍ��o\g8tt��| e���Rw����S�0�X4w�Ų�L+���j�]�YKK#�Qt��K��a����|�d�eGX[��<��)C�Z�X��.f�U�>j"YQ��5B����=�����<�W�̴����'k�`o��BFLʧg�=��X7$s?��I��-f�A�Z��4��N+�ElH��hϭ�g( (�j���d�$X��{ Ⴘ���&!)T��!�)u�b.]�������񻃶f�	�ܧ�KYr�g%���3��>�,�P�V�6֠��z��@z+���)
�����ヤx��2�m�Kc)o�4HE�陕}�"%�V����p3�C��-K����6�N8�����	U"��ȸ{�zڇ�o1��w���i���g9��v*W�E��Q�ŌZy��~R�%�T�u^��x�)r~Y@g��h�ǁ��
���3��*��E�l�5K�E��x!��Jß^;����؞(S��f��M�s띋偃2� ��>�Ƈ�tw7�Y[Xlt&P
�׸ۼ���������6vij��5T����NH�gj'�d�:9��Q�k���a�ͧ�B�����OE#�UX�jaE�J�+�mm��7Շjc����8(��gh��	[u��8f��V"��^0ؚY��#�[<�v��wܐ�j�o��� ����a�!��.�w�Uw�!��\"�IwJ?��p\��s�u�1�v����:")�'��� x����w�9T��[��N⧂�K�^�%�A��՞��.̈:,�P����������IY:m��;lɖ|�0�� �(���(�O�4\�=)�o�q!i3��zD�J�ZY>�-e�וWl.�Τmd:ir+뿆٫b�~-�F޲�{�	Ys?]�a���!.��=E���Sa�WPB2jMM�H���CCe6�@B3�Q���sr�ARr�w��[�hd� :�z,��9���a:ry�����F��k4�%�FW��^�ֺ��$}7R��m>�Kv"^30�x[�8�SX��҉$��.��+Pl4y����������l��V�U����������;�B�r�� "��=�,���=E2��E������!u�Z)#���F'ؚ����\�4v ��5:0�k���A����.Y�`���?Z�	��6����Ad�U�{X��y�QSM�2A�`��t&;:���0UT�˽���4%�_^���Lc-��TEn�/`����,QL���kc9A�=F8_2	��~5�*8O�
��d﵏�mu��=�u�gN�'��z��ԑ � ��.%��ޑX$*�咽y�xĬC᫵�w����t�k�8�JF)*Z�d��M���
�fҧ�r�f�O�ਖ਼�y��܇;�0�C�5�8���Z.�>3IV0���j�c� ����~yH���t�.#ZF`�Z����w�2 Ͽk,o�-�A�� G�1b(d8��!Y�/|���I��s�2��A�⥁zV��ڃ�3`c�}DC��Wm�{�>í���I3��k�C#r�3J��>i�E�1,&ν��|�f4�!v����J$�Za W��#>-���u��6>w� �/�rBiYd�v���ү�謞7��N�:"�q�������w��%	�[�v��(�(�%�XȾ�k��Da�{�U��p��RsΦ�N�C��\��p��oU�K��U���#H��-SY�lݐ�i�l�F)�*�ј���mv�%�#.�p��'���P=O�אTW��hQ�/&�2[�h�텸x�E��õ �$2� �M]$�*fnЩ��b�� Kv9=<.�ˁ�������s��y�A�OWKN�A���71?�K�$!!t��M�
��:056����KcB��CH������tXp�U�<pq�5��.<�$��s^��(�Ya�H~W��-*�
���g�mɬ���3��gz�H&�:G�IQU�6ܭ�o��\}�}�{߆�G���H�wU�
4��$p������X����o�Ȱ[`-9��k�m�2z90n���f��������H�
�Hw����$�έgʶ�ņw��&�vbI�*WN�FE_	y@`W�g��4�Xq�n�H����j��u|p�5J�&�x�E��~x�ޱ�	�Lᇰݱ���s���{�)���+�����Da�X�2-g�ט#�>�r�]�P��a��)�׃���s���P��`�K4'k#��/���$��GҲ$6�7���^�;I��)q;���~z��}��H.8��B�"�"�F2m^�̃$�����jt���k�md��uH�,=e�����U��= ��OR���B�,�w�~�������}f`�e�m6e����GԠu@�ɷ��Wn��[؇KHI�>>Z��[i��3��ymt�>�^�*ݙ�/r`,ShRlm]�垫-+��9m{�}����3�>�a蠽}�:x@���2�v����х� `F�+S��j�~dC����9`��O��$˗ze���)����$��9d��\`.���-QE�����4���Lg�g�I����Ą[�Q6�k ��s�1��W��Y:i@�4c7Q~j��HE��|��C/��IE�>`z�>!_p��Y�K��ȓ-��J��<x�f�M^R��|&�oڊ���ˑ�3�H�E3)��X�}�H:Wgh��(K�V�U��KX� ,��׻d7_~��\���Ibɶ��x5�+��m������6�6�s�`a�x?��%��FA��~\���w���[ó����4�ˣ�%eͩA�S��\>�	^�$w������?���l��X�x;��H�AӚ��iCE����Q/����q)3'�e��y\�s�؄U"��*����xy�?b�|;,�<��jt��+�Wj������uͩ�iDd.��I�	~uy����_D�Lb*.��J1�TN�-yU��|l��Ǚrrl�)��fI�* �\��})�Ч��+�!����fo�/�I~\I�=%<�.g7�r7V���7n���ڹQ)\�:]Z���$��<��GU�&9U��V�ÃLf�=�b8��ǴcKj�hW'���� Cn3��*��I�I�
#���1u�>��nttE��q�����(���<���� ���D&��L��,��Uy+�����~),�,�����TcK)�bs�/�!v�*�<Ųh��ܟ��-��M��9���%���R��a�7�1�����u�g �8���z�8�u7��1��".������*^�b]p���ƥ2� �:�2I�ف�������,��9<��>�#��l���"U]����d�Rz��� !DE�F�~x`W�C�+JY(N�85������K~��$����c�_:"Da�]����x�(��B/C�uK��;���v������?���W�X$�NɊ��0mi�P�6膪��s���3�����nA�'X�fX6#n8�e��b��S|�鑀]"E	���#@��D6�] ꝲ�1m�+�@i���Zp3H;�s�a����V�-�s��6;��N��x�r��Fۏ���;ǩ{2d�"[ :
?���	%� ���<���i����e˟�m�|�>l�����;�
���FPIp�qۥ~���? �y>���g+&��f�zl������!g�j鯱_M4��&W>T��f#�s����C�J�ӝ-�k��f��;=ɠ~d m	��5�B��T9_����	�=."!*Wb	v�j�8@�W��!����c��ː%���o������ ���(C~�Q=��R�5o�L,ƿ���y����q�t���Χ�� �y*�p|	0\@��y��(C��9_(�X{��@w�p��We�5�^���"��61�'q={�xRS��=��ͷ8�ƒ'��s���rɷ:O-� t9���wp�fJ�\%%�pM�ٽ`+���{f�7��1�2�m��+Љ�5��?�����ɟ��x���Q"`�P̔Fm�Ijj�rq	�|Ц#�O����ʝ��w����D���(�?��yY��Ο3]-4��)z	P��y�ˊ�a�#��1�E�]��F:#���Jssp'�e���R����w�e��F��GR%�S��՟	&x��K]ڼ�U]���p�V=4{p>�6�1��m	��z�D�!Z��P��u����^#�,�.!T��*��@�H��=ms��v+�7���q����t���ӚFJɱ_7�R���P_��h~� CE��&ڳuݥ#lOl����n�w��ޑ� ��|���u�Ax��q4�����.2:}���%��Z��G�
Y���C㕸�^�La3�"����/�Y�7����X�� ��շܠ�%v�.�t��V,�qp�9`�_;c&�����M���+ �[�ʉ!h/|�#�mx����ƫ�X�qfoj�
+���ڕP���}�^	گ���\ �a�}wA�VL�������*�5�ez�\� nTQw�^��(�{�5BGM+��B���B�n�In��z��J��A�%����5 .��mjd�\v2���YD�RlK�#=���I@�F �I%i�!���vB|�6)u*��	AT�	��:����=�0����䆉�E�Q�@���8�e���&���9��m�Z]���t���V�ҿ�^�0L*�`��B�t�[�L�&�����Ƕ8`����ID,�[�FUR��
|J#w�d#H}�:i���J]<�ً���}��:��糾
��u�j�3�O�����$��m ���ܠ��P�`祝���Y7��i!:��!�ٜ�+8K`w��1	�|�]eY:�5%唵Y�
H>!�rLE�3�@ܢ9:�k��i��@�rF�-.���3٥���
Zz����.8����*��$��j�K'���z�&����k��Z���0fv�4 \�'�	�u7�iT�"�b��n�em�~PKI �&v��E���q >�>h1o�I�^�) �D絴�Q(J���Z�n�V� M�^V�3K1T��� ���;����)��A�i6�2}�a�P<b �VW!ȓ�Ds���� ߅��n�&�g�uP���4��w�_������I�.�����X�[x.s��C� �i)wf:��V�őlS��ʾ��,�)o7�ՂC+���:./�ݟ�A~���Y���i���aO�X�^E6|��i{ �}�l�)�l(��.u�0��S�����0���'P܆�c�e���ڪG	+F�I�& ��nۅ[�%�Ӛ�D�.��w��) a�Y	�@��=�<��r���@V'-�Ӹ�ϔ�P��\��Y$��=e8���P^��:`�H�q��0 T�U9�y�q����;kAՉ��6徉\��7Ҷ샢5��X�"���]�-m=32fPe�ŕ���KV�
��f�0lV�R��n�%�`C^�Q9����%�p�\�A�����e���f��N"����yG�#|uMaoG��LI�N������r�����ߚ:��|
�c-�UAJ�(���4��+F����)���p��U�g��x3� �+��Z�����{��]��P��ao;G�&r�mj[��r3+��kPp�	� ��
_u�ⅆ�p�B���כ
.��	��2�y�%}8��W��dg2�m�Du�Lx=<'.�	��f�^sZ�̸���w��(�w��)Q�Q�o�|?F�N�|[j'*��evI��:�Z�:��H�5�S(��sC �?&,�K�֑�
/��Ӓ4�^�.R^��̧o�8P������������~�lAk%sB������F@�J��!`E��A�N�J���I��|��Es�v���'��H�+�I���%���^Myo�� � ��%W�w�)]����~�z!��o PAZ��8�TK�F�S(Ú�쪗�����k�G�yU��ҏE)��<�Ɣ埽��o�/j|��R���:|v��+c׭:�'��S��K�5��P��Eٷ�ᓤ��\������<!,�S���d�H���������h��7��
U�H?����_	19�j���i�����#E�������v1���N��.�uM��ͅ�
F�YɌ�?�à,��āV!tX�����[:=1�Z�fZ����*^#�vc��,9P���ф`��fp���u0%ޱ*�l&h,�L�ȈJ/u�����SY��P�tҍ5���f�j�mc����"y����}iM#\��W��}#L�@�XFՍ4d[jtUž�[D.�de�7�+������R��E��#�)j�7�>O�WL�:��D�ϙ�S%ORv��#�!P�i�FR�νׄR��F8�%8U�mR��zL�(qF之�6�C%~C������P�(���80�TT�-��GҸ��	�;�xZ����ݙ�rdµCe͚�e��6N�6�=������:b*��������"����i���P��y��^`j�oj�S����$C�ˡ�杢���K�aQ�`iﰴ�y��,z�M�.2�!B`��J�mmK��]�$s�3F��oV����y�j�Bp��۫�g���T�J���0|��*��eL�[#
��Pl�':��
U"Tи�!���d.0H��Pݰ���<��l�~�"$dՇ���u�1����ߨl�B�'.IR�������/T*���
��$�w�`TGf���|��L���#��W�I+�c�J'�A���	a*��oj~<�U����~z�6ZE���a��0�0����Z����(#�##�/5U_��$�C�~|�^� ����x�}7Y7φ	0����E��j>I"6��L��؍����r'�l.�w����Ќ����0�6�0����a|��������jem+��1�[�n�ѵ�S�㆞+L]�V�'!ked�	�a1q�P����W�i�AǾ �iR�U,��#y�B��W�1X"0�K�q4-�(�/M{P{�Df��hCGK�%��,�[�R�?���Y��/�,�GΡ3~8^��U��7����Y@�R�R,�Ɓj�-��n�����7�DES�		�e[ؗ��	�g��9q���?BF$���?%�rz���
n/I��ߏNz�jf\�Xز���m5�f�-S�l;�G�x�T����a��I�Rh��ۛ�1Ol!O[��V��O9�J��.ćY�r�EF��_���=���s�ܮ�5�6���e�<*��e�����y�e�¬��v�w4���E%wD��hrd:�w��%��y�/�jw�b��1<��ՖF�P��;��ǎ���ە���+V�^�;LC�����v��53o/M���4�{�J�%ZTL;@��O��nWi�R\���_��p��4T{�`�>�p�����ʅdf�{�7/:gcg�լX8v��� ��FN���̀��yxTS����6lY��ٞ�-G�ޚֈg�0���0߹�aP�����f��_�%ɋ�:�0�X��j_�a�����P��	��-a������5++���W/��}n�~���@��?�.iHVe��6�\N���Mл�Ŝ}v�὾��BFqb7�F3$֕8{K����� ��/v]���g�h׮��y��U��ح��0֦�^�4�c��Y羇Ȼ9�H�^)i8eB�4��W��(M��}��uVN�`C��m�h�~�W�|�g��'�lUqy�k��f�-�~�k�f�l�K�«1��~��/֙�f�r���E9���Q��ɲB(�ђ��w���R��~VM<���R���t2��V�PN���K�*_z��޽����{�G��q�[��A*��lQK�HVV,�7�I%A(2;�1�p�9H��ŌP��Ң��'y�S�ķ�n�]�8C��߷��)��K�i�A�lT�� �/�~�ߓ�Mu�ڈ,���Z/��E��?�n�bS`��$���q����а����x 'O%�Ս9Z��m���_�u��R����,��<�v��&_�Q����<�#�ҔW�jy��qT2����0P%P�i`S��.�۲1Z<k�x��f_հμ��2������v�*���_F���f�D.����@H0��=�y�v%�h�����Q��T0ؤ�n�� '�{@�t��]{��C/u�tE��L�l:fI����^�X9j`��e�#
�֋�����h
ƃD Ժ��o�{,�(zĝ{x� U��U��oc)O�sS�/�5b��&����0(2寳�eE�ܩ\<�c�1��lK᜞��܌IVg5lPkZ�|�qڙ;eƂf�v��E�0��@1-]�h�B���q����̆㟀V�B�H7{����Lb�JY5/,`	^